----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/17/2022 04:16:05 PM
-- Design Name: 
-- Module Name: phaser_datapath_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

use STD.textio.all;
use ieee.std_logic_textio.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity phaser_datapath_tb is
--  Port ( );
end phaser_datapath_tb;

architecture Behavioral of phaser_datapath_tb is
    constant half_period: time := 10ns;
    signal on_in_s : STD_LOGIC;
    signal clk :  STD_LOGIC := '0';
    signal input_in_s : STD_LOGIC_VECTOR (15 downto 0) := x"0000";
    signal output_out_s : SIGNED(15 downto 0);
    signal reset : std_logic;
    signal out_valid: std_logic;
    
    signal input_from_file_s: STD_LOGIC_VECTOR (15 downto 0);
    type audio_type is array (441343 downto 0) of std_logic_vector(15 downto 0);
    
    signal AUDIO : audio_type :=(
    "1111111111110111",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010011",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000001001",
    "0000000000001110",
    "0000000000010011",
    "0000000000010110",
    "0000000000011001",
    "0000000000011001",
    "0000000000010111",
    "0000000000010110",
    "0000000000010011",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001111",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010011",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000001111",
    "0000000000001100",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000010",
    "1111111111111100",
    "1111111111110111",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110111",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101101",
    "1111111111101010",
    "1111111111100111",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001110",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001100",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001100",
    "0000000000001001",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000000",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000100",
    "0000000000000111",
    "0000000000001100",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001001",
    "0000000000000101",
    "1111111111111110",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "0000000000000100",
    "0000000000001010",
    "0000000000001111",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010001",
    "0000000000001100",
    "0000000000000101",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000000111",
    "0000000000000000",
    "1111111111111001",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101010",
    "1111111111101100",
    "1111111111101101",
    "1111111111110001",
    "1111111111110110",
    "1111111111111001",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001100",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000010",
    "1111111111111011",
    "1111111111110111",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110111",
    "1111111111111011",
    "0000000000000010",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000100",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111110",
    "0000000000000101",
    "0000000000001010",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001001",
    "0000000000000100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000101",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111100",
    "0000000000000010",
    "0000000000001001",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001001",
    "0000000000000101",
    "0000000000000000",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000100",
    "1111111111111110",
    "1111111111111001",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "0000000000000000",
    "0000000000000101",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111011",
    "0000000000000010",
    "0000000000000111",
    "0000000000001110",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010001",
    "0000000000001100",
    "0000000000000111",
    "0000000000000010",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111011",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101111",
    "1111111111110010",
    "1111111111110111",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111101111",
    "1111111111101010",
    "1111111111100111",
    "1111111111100100",
    "1111111111100010",
    "1111111111100100",
    "1111111111100101",
    "1111111111101001",
    "1111111111101101",
    "1111111111110010",
    "1111111111111001",
    "1111111111111110",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000000101",
    "1111111111111100",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000000",
    "1111111111111011",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101101",
    "1111111111101101",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001010",
    "0000000000000111",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010100",
    "0000000000010011",
    "0000000000010001",
    "0000000000001110",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000000111",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "0000000000000000",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111100",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111110110",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001010",
    "0000000000000101",
    "1111111111111110",
    "1111111111111001",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111001",
    "1111111111110100",
    "1111111111101111",
    "1111111111101100",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111110001",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000001001",
    "0000000000001100",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "0000000000000000",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001100",
    "0000000000001111",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010011",
    "0000000000001111",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111110",
    "0000000000000100",
    "0000000000001001",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001110",
    "0000000000010011",
    "0000000000010111",
    "0000000000011100",
    "0000000000100001",
    "0000000000100101",
    "0000000000100110",
    "0000000000100101",
    "0000000000100000",
    "0000000000010111",
    "0000000000001110",
    "0000000000000010",
    "1111111111110010",
    "1111111111100111",
    "1111111111011101",
    "1111111111010111",
    "1111111111010010",
    "1111111111010000",
    "1111111111010010",
    "1111111111010111",
    "1111111111011101",
    "1111111111100101",
    "1111111111101111",
    "1111111111110111",
    "0000000000000010",
    "0000000000001001",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001100",
    "0000000000000111",
    "0000000000000010",
    "1111111111111011",
    "1111111111110110",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111110001",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000000",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000000",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001110",
    "0000000000001100",
    "0000000000001010",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000001001",
    "0000000000001010",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000100",
    "0000000000001010",
    "0000000000010001",
    "0000000000011001",
    "0000000000100000",
    "0000000000101000",
    "0000000000101110",
    "0000000000110010",
    "0000000000110101",
    "0000000000110011",
    "0000000000110000",
    "0000000000101000",
    "0000000000011100",
    "0000000000001111",
    "1111111111111110",
    "1111111111101111",
    "1111111111100010",
    "1111111111010111",
    "1111111111010010",
    "1111111111010000",
    "1111111111010010",
    "1111111111011010",
    "1111111111100101",
    "1111111111110010",
    "0000000000000010",
    "0000000000001111",
    "0000000000011001",
    "0000000000100001",
    "0000000000100101",
    "0000000000100110",
    "0000000000100101",
    "0000000000100001",
    "0000000000011100",
    "0000000000010111",
    "0000000000010001",
    "0000000000001100",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000000",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000001110",
    "0000000000010100",
    "0000000000011001",
    "0000000000100000",
    "0000000000100011",
    "0000000000100101",
    "0000000000100101",
    "0000000000100001",
    "0000000000011100",
    "0000000000010011",
    "0000000000000111",
    "1111111111110111",
    "1111111111101010",
    "1111111111011111",
    "1111111111010111",
    "1111111111010010",
    "1111111111010000",
    "1111111111010000",
    "1111111111010101",
    "1111111111011011",
    "1111111111100101",
    "1111111111101101",
    "1111111111110111",
    "0000000000000010",
    "0000000000001001",
    "0000000000001110",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001001",
    "0000000000000101",
    "0000000000000000",
    "1111111111111001",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101010",
    "1111111111101010",
    "1111111111101100",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110110",
    "1111111111110111",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "0000000000000000",
    "0000000000000101",
    "0000000000001010",
    "0000000000001110",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010011",
    "0000000000001111",
    "0000000000001100",
    "0000000000000111",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111110",
    "0000000000000111",
    "0000000000001110",
    "0000000000010100",
    "0000000000011011",
    "0000000000100001",
    "0000000000100110",
    "0000000000101011",
    "0000000000101011",
    "0000000000101000",
    "0000000000100001",
    "0000000000010111",
    "0000000000001010",
    "1111111111111011",
    "1111111111101111",
    "1111111111100100",
    "1111111111011101",
    "1111111111011011",
    "1111111111011011",
    "1111111111011101",
    "1111111111100010",
    "1111111111101001",
    "1111111111101111",
    "1111111111110111",
    "0000000000000000",
    "0000000000000111",
    "0000000000001110",
    "0000000000010001",
    "0000000000010100",
    "0000000000010110",
    "0000000000010110",
    "0000000000010110",
    "0000000000010110",
    "0000000000010100",
    "0000000000010001",
    "0000000000001110",
    "0000000000001001",
    "0000000000000100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000101",
    "0000000000001001",
    "0000000000001110",
    "0000000000010001",
    "0000000000010100",
    "0000000000010111",
    "0000000000011011",
    "0000000000011110",
    "0000000000100000",
    "0000000000100011",
    "0000000000100101",
    "0000000000100011",
    "0000000000100000",
    "0000000000011001",
    "0000000000010011",
    "0000000000001100",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000001010",
    "0000000000010001",
    "0000000000011001",
    "0000000000100011",
    "0000000000101011",
    "0000000000110011",
    "0000000000111010",
    "0000000000111101",
    "0000000000111111",
    "0000000000111011",
    "0000000000110111",
    "0000000000110000",
    "0000000000100101",
    "0000000000011001",
    "0000000000001110",
    "0000000000000000",
    "1111111111110100",
    "1111111111101100",
    "1111111111100101",
    "1111111111100010",
    "1111111111100100",
    "1111111111100111",
    "1111111111101101",
    "1111111111110100",
    "1111111111111100",
    "0000000000000111",
    "0000000000001110",
    "0000000000010100",
    "0000000000011001",
    "0000000000011100",
    "0000000000011100",
    "0000000000011011",
    "0000000000011001",
    "0000000000010110",
    "0000000000010011",
    "0000000000001110",
    "0000000000001001",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "0000000000000100",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "0000000000000100",
    "0000000000001001",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110110",
    "1111111111110001",
    "1111111111101010",
    "1111111111100101",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100101",
    "1111111111100111",
    "1111111111101100",
    "1111111111110001",
    "1111111111110110",
    "0000000000000000",
    "0000000000001100",
    "0000000000010111",
    "0000000000100001",
    "0000000000101001",
    "0000000000101110",
    "0000000000101110",
    "0000000000101101",
    "0000000000101000",
    "0000000000100101",
    "0000000000100000",
    "0000000000011110",
    "0000000000011011",
    "0000000000011001",
    "0000000000011001",
    "0000000000011011",
    "0000000000011110",
    "0000000000100101",
    "0000000000101001",
    "0000000000110000",
    "0000000000110011",
    "0000000000110011",
    "0000000000101110",
    "0000000000100101",
    "0000000000010110",
    "0000000000000010",
    "1111111111101100",
    "1111111111010101",
    "1111111111000001",
    "1111111110101111",
    "1111111110100010",
    "1111111110011010",
    "1111111110010111",
    "1111111110011000",
    "1111111110011101",
    "1111111110100101",
    "1111111110110001",
    "1111111110111100",
    "1111111111001011",
    "1111111111011010",
    "1111111111100111",
    "1111111111110001",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101101",
    "1111111111101001",
    "1111111111100100",
    "1111111111011111",
    "1111111111011011",
    "1111111111011000",
    "1111111111010111",
    "1111111111011010",
    "1111111111011101",
    "1111111111100010",
    "1111111111100111",
    "1111111111101100",
    "1111111111101111",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100101",
    "1111111111100101",
    "1111111111100101",
    "1111111111100111",
    "1111111111101001",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001100",
    "0000000000010001",
    "0000000000010110",
    "0000000000011001",
    "0000000000011100",
    "0000000000011110",
    "0000000000011110",
    "0000000000011011",
    "0000000000011001",
    "0000000000010100",
    "0000000000010011",
    "0000000000010011",
    "0000000000010100",
    "0000000000010111",
    "0000000000011001",
    "0000000000011011",
    "0000000000011011",
    "0000000000010111",
    "0000000000010100",
    "0000000000010011",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010110",
    "0000000000011001",
    "0000000000100000",
    "0000000000100101",
    "0000000000101011",
    "0000000000110000",
    "0000000000110010",
    "0000000000110011",
    "0000000000110000",
    "0000000000101011",
    "0000000000100101",
    "0000000000011100",
    "0000000000010011",
    "0000000000001010",
    "0000000000000010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "0000000000000000",
    "0000000000000111",
    "0000000000001010",
    "0000000000001111",
    "0000000000010100",
    "0000000000011001",
    "0000000000011100",
    "0000000000100000",
    "0000000000100011",
    "0000000000100101",
    "0000000000100110",
    "0000000000100110",
    "0000000000100101",
    "0000000000100011",
    "0000000000011110",
    "0000000000011001",
    "0000000000010011",
    "0000000000001110",
    "0000000000001010",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "0000000000000010",
    "0000000000000111",
    "0000000000001100",
    "0000000000001111",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010100",
    "0000000000010100",
    "0000000000010011",
    "0000000000010001",
    "0000000000001110",
    "0000000000001100",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000101",
    "0000000000000000",
    "1111111111111011",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101100",
    "1111111111101101",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110010",
    "1111111111101101",
    "1111111111101001",
    "1111111111100101",
    "1111111111100100",
    "1111111111100111",
    "1111111111101010",
    "1111111111110010",
    "1111111111111100",
    "0000000000001010",
    "0000000000010100",
    "0000000000100000",
    "0000000000101000",
    "0000000000101110",
    "0000000000110000",
    "0000000000101110",
    "0000000000101000",
    "0000000000100000",
    "0000000000010011",
    "0000000000000101",
    "1111111111110110",
    "1111111111101010",
    "1111111111100010",
    "1111111111011011",
    "1111111111010111",
    "1111111111010101",
    "1111111111010101",
    "1111111111011000",
    "1111111111011101",
    "1111111111100101",
    "1111111111101101",
    "1111111111110111",
    "0000000000000010",
    "0000000000001001",
    "0000000000001111",
    "0000000000010011",
    "0000000000010011",
    "0000000000010001",
    "0000000000001100",
    "0000000000000111",
    "1111111111111100",
    "1111111111110110",
    "1111111111101101",
    "1111111111101001",
    "1111111111100101",
    "1111111111100100",
    "1111111111100101",
    "1111111111101001",
    "1111111111101111",
    "1111111111110111",
    "0000000000000010",
    "0000000000001010",
    "0000000000001111",
    "0000000000010011",
    "0000000000001111",
    "0000000000001010",
    "1111111111111110",
    "1111111111110010",
    "1111111111100111",
    "1111111111011011",
    "1111111111010101",
    "1111111111010010",
    "1111111111010010",
    "1111111111010111",
    "1111111111011101",
    "1111111111100111",
    "1111111111101111",
    "1111111111111001",
    "0000000000000100",
    "0000000000001100",
    "0000000000010100",
    "0000000000011100",
    "0000000000100101",
    "0000000000101001",
    "0000000000101101",
    "0000000000110000",
    "0000000000110000",
    "0000000000110010",
    "0000000000110011",
    "0000000000110111",
    "0000000000111000",
    "0000000000111010",
    "0000000000111101",
    "0000000000111101",
    "0000000000111101",
    "0000000000111011",
    "0000000000111010",
    "0000000000110111",
    "0000000000110010",
    "0000000000101110",
    "0000000000101000",
    "0000000000100001",
    "0000000000010111",
    "0000000000001110",
    "0000000000000010",
    "1111111111110100",
    "1111111111101001",
    "1111111111011101",
    "1111111111010101",
    "1111111111010000",
    "1111111111001011",
    "1111111111001001",
    "1111111111001011",
    "1111111111001101",
    "1111111111010000",
    "1111111111010011",
    "1111111111010111",
    "1111111111011011",
    "1111111111011111",
    "1111111111100000",
    "1111111111100100",
    "1111111111100101",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100111",
    "1111111111100101",
    "1111111111100101",
    "1111111111100101",
    "1111111111100101",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100101",
    "1111111111100100",
    "1111111111100100",
    "1111111111100101",
    "1111111111100111",
    "1111111111101010",
    "1111111111101100",
    "1111111111101100",
    "1111111111101010",
    "1111111111100111",
    "1111111111100010",
    "1111111111011101",
    "1111111111011000",
    "1111111111010101",
    "1111111111010101",
    "1111111111010101",
    "1111111111011010",
    "1111111111100000",
    "1111111111100111",
    "1111111111110001",
    "1111111111111011",
    "0000000000000111",
    "0000000000001111",
    "0000000000010111",
    "0000000000011100",
    "0000000000100000",
    "0000000000100001",
    "0000000000100000",
    "0000000000011011",
    "0000000000010100",
    "0000000000001001",
    "1111111111111001",
    "1111111111101100",
    "1111111111011011",
    "1111111111001110",
    "1111111111000011",
    "1111111110111001",
    "1111111110110110",
    "1111111110110110",
    "1111111110111011",
    "1111111111000011",
    "1111111111001110",
    "1111111111011011",
    "1111111111101010",
    "1111111111111001",
    "0000000000000111",
    "0000000000010011",
    "0000000000011011",
    "0000000000011110",
    "0000000000011100",
    "0000000000011001",
    "0000000000010011",
    "0000000000001110",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000000111",
    "0000000000000100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "0000000000000010",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010011",
    "0000000000010100",
    "0000000000010111",
    "0000000000011011",
    "0000000000011110",
    "0000000000100001",
    "0000000000100011",
    "0000000000100101",
    "0000000000100101",
    "0000000000100101",
    "0000000000100101",
    "0000000000100101",
    "0000000000100110",
    "0000000000101000",
    "0000000000101000",
    "0000000000100110",
    "0000000000100101",
    "0000000000100001",
    "0000000000100000",
    "0000000000011100",
    "0000000000011011",
    "0000000000011011",
    "0000000000011001",
    "0000000000010110",
    "0000000000010011",
    "0000000000010001",
    "0000000000001110",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010011",
    "0000000000010100",
    "0000000000010110",
    "0000000000010110",
    "0000000000010110",
    "0000000000010110",
    "0000000000010110",
    "0000000000010111",
    "0000000000011001",
    "0000000000011001",
    "0000000000011100",
    "0000000000011100",
    "0000000000011100",
    "0000000000011100",
    "0000000000011011",
    "0000000000010111",
    "0000000000010100",
    "0000000000010001",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000010001",
    "0000000000010110",
    "0000000000011110",
    "0000000000100110",
    "0000000000101110",
    "0000000000110111",
    "0000000000111010",
    "0000000000111011",
    "0000000000111000",
    "0000000000110011",
    "0000000000101001",
    "0000000000011110",
    "0000000000010011",
    "0000000000000111",
    "1111111111111011",
    "1111111111110010",
    "1111111111101101",
    "1111111111101010",
    "1111111111101100",
    "1111111111101101",
    "1111111111110010",
    "1111111111111001",
    "0000000000000100",
    "0000000000001100",
    "0000000000010011",
    "0000000000011001",
    "0000000000011110",
    "0000000000100000",
    "0000000000100001",
    "0000000000100001",
    "0000000000100000",
    "0000000000011110",
    "0000000000011100",
    "0000000000011100",
    "0000000000011011",
    "0000000000010111",
    "0000000000010100",
    "0000000000010001",
    "0000000000001100",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111101001",
    "1111111111101001",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101101",
    "1111111111110010",
    "1111111111110111",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101100",
    "1111111111101101",
    "1111111111110010",
    "1111111111111001",
    "0000000000000100",
    "0000000000001100",
    "0000000000010011",
    "0000000000011001",
    "0000000000011100",
    "0000000000011100",
    "0000000000011001",
    "0000000000010011",
    "0000000000001001",
    "1111111111111011",
    "1111111111101111",
    "1111111111100101",
    "1111111111011011",
    "1111111111010101",
    "1111111111010010",
    "1111111111010000",
    "1111111111010000",
    "1111111111010000",
    "1111111111010000",
    "1111111111010010",
    "1111111111010011",
    "1111111111010111",
    "1111111111011011",
    "1111111111100010",
    "1111111111101001",
    "1111111111110001",
    "1111111111111001",
    "1111111111111110",
    "0000000000000100",
    "0000000000000101",
    "0000000000000101",
    "0000000000000101",
    "0000000000000100",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001100",
    "0000000000010011",
    "0000000000011100",
    "0000000000101001",
    "0000000000110111",
    "0000000001000100",
    "0000000001010001",
    "0000000001011011",
    "0000000001100000",
    "0000000001011110",
    "0000000001010110",
    "0000000001001001",
    "0000000000110111",
    "0000000000100011",
    "0000000000001110",
    "1111111111110110",
    "1111111111100010",
    "1111111111010000",
    "1111111111000001",
    "1111111110110110",
    "1111111110101100",
    "1111111110100111",
    "1111111110100101",
    "1111111110101001",
    "1111111110101100",
    "1111111110110010",
    "1111111110111011",
    "1111111111000011",
    "1111111111001011",
    "1111111111010101",
    "1111111111011011",
    "1111111111100010",
    "1111111111100111",
    "1111111111100111",
    "1111111111100111",
    "1111111111100101",
    "1111111111100010",
    "1111111111011111",
    "1111111111011011",
    "1111111111011010",
    "1111111111011000",
    "1111111111011010",
    "1111111111011011",
    "1111111111011111",
    "1111111111100000",
    "1111111111100101",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100100",
    "1111111111100000",
    "1111111111011101",
    "1111111111011010",
    "1111111111010111",
    "1111111111010101",
    "1111111111010011",
    "1111111111010011",
    "1111111111010101",
    "1111111111010101",
    "1111111111011000",
    "1111111111011010",
    "1111111111011010",
    "1111111111011011",
    "1111111111011011",
    "1111111111011011",
    "1111111111011011",
    "1111111111011011",
    "1111111111011101",
    "1111111111011111",
    "1111111111100000",
    "1111111111100010",
    "1111111111100101",
    "1111111111100111",
    "1111111111101001",
    "1111111111101001",
    "1111111111101001",
    "1111111111101001",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101100",
    "1111111111101101",
    "1111111111110010",
    "1111111111110111",
    "1111111111111011",
    "0000000000000010",
    "0000000000000101",
    "0000000000001001",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010100",
    "0000000000010111",
    "0000000000011001",
    "0000000000011001",
    "0000000000011011",
    "0000000000011100",
    "0000000000011100",
    "0000000000011100",
    "0000000000011100",
    "0000000000011001",
    "0000000000010110",
    "0000000000010011",
    "0000000000001111",
    "0000000000001100",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001010",
    "0000000000001100",
    "0000000000001110",
    "0000000000001111",
    "0000000000001111",
    "0000000000010001",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010110",
    "0000000000011001",
    "0000000000011100",
    "0000000000100001",
    "0000000000101000",
    "0000000000101011",
    "0000000000101110",
    "0000000000110000",
    "0000000000101110",
    "0000000000101011",
    "0000000000100110",
    "0000000000100000",
    "0000000000011011",
    "0000000000011001",
    "0000000000011001",
    "0000000000011011",
    "0000000000100001",
    "0000000000101001",
    "0000000000110010",
    "0000000000111101",
    "0000000001000111",
    "0000000001010001",
    "0000000001010110",
    "0000000001011001",
    "0000000001010111",
    "0000000001010010",
    "0000000001001001",
    "0000000000111111",
    "0000000000110010",
    "0000000000100110",
    "0000000000011100",
    "0000000000010011",
    "0000000000001010",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001100",
    "0000000000010011",
    "0000000000011001",
    "0000000000100000",
    "0000000000100110",
    "0000000000101101",
    "0000000000110010",
    "0000000000110101",
    "0000000000110111",
    "0000000000110111",
    "0000000000110011",
    "0000000000110000",
    "0000000000101011",
    "0000000000100110",
    "0000000000100011",
    "0000000000100000",
    "0000000000011110",
    "0000000000011100",
    "0000000000011100",
    "0000000000100000",
    "0000000000100001",
    "0000000000100101",
    "0000000000100110",
    "0000000000101000",
    "0000000000100110",
    "0000000000100011",
    "0000000000100000",
    "0000000000011011",
    "0000000000010111",
    "0000000000010110",
    "0000000000010110",
    "0000000000010111",
    "0000000000010111",
    "0000000000010111",
    "0000000000010110",
    "0000000000010100",
    "0000000000010001",
    "0000000000001111",
    "0000000000001110",
    "0000000000001100",
    "0000000000001100",
    "0000000000001100",
    "0000000000001110",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010100",
    "0000000000010011",
    "0000000000001111",
    "0000000000001110",
    "0000000000001001",
    "0000000000000101",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101100",
    "1111111111100101",
    "1111111111011111",
    "1111111111011011",
    "1111111111011010",
    "1111111111011010",
    "1111111111011101",
    "1111111111100010",
    "1111111111100111",
    "1111111111101101",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110001",
    "1111111111101010",
    "1111111111100100",
    "1111111111011101",
    "1111111111011010",
    "1111111111011000",
    "1111111111011000",
    "1111111111011011",
    "1111111111100010",
    "1111111111101010",
    "1111111111110100",
    "1111111111111110",
    "0000000000001010",
    "0000000000010001",
    "0000000000010110",
    "0000000000010110",
    "0000000000010100",
    "0000000000010001",
    "0000000000001010",
    "0000000000000100",
    "1111111111111001",
    "1111111111110001",
    "1111111111101001",
    "1111111111100000",
    "1111111111011000",
    "1111111111010011",
    "1111111111010000",
    "1111111111001101",
    "1111111111001110",
    "1111111111010000",
    "1111111111010010",
    "1111111111010101",
    "1111111111011000",
    "1111111111011011",
    "1111111111011111",
    "1111111111100000",
    "1111111111100100",
    "1111111111100111",
    "1111111111101100",
    "1111111111101111",
    "1111111111110100",
    "1111111111111011",
    "0000000000000100",
    "0000000000001001",
    "0000000000001110",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001100",
    "0000000000000111",
    "0000000000000010",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111101111",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100101",
    "1111111111100010",
    "1111111111100000",
    "1111111111011101",
    "1111111111011011",
    "1111111111011000",
    "1111111111010111",
    "1111111111010101",
    "1111111111010011",
    "1111111111010010",
    "1111111111010010",
    "1111111111010011",
    "1111111111010011",
    "1111111111010101",
    "1111111111011000",
    "1111111111011101",
    "1111111111100100",
    "1111111111101100",
    "1111111111110100",
    "1111111111111110",
    "0000000000001001",
    "0000000000010011",
    "0000000000011100",
    "0000000000100101",
    "0000000000101101",
    "0000000000110101",
    "0000000000111000",
    "0000000000111011",
    "0000000000111011",
    "0000000000111010",
    "0000000000110111",
    "0000000000110000",
    "0000000000101001",
    "0000000000100011",
    "0000000000011100",
    "0000000000010100",
    "0000000000001110",
    "0000000000000101",
    "1111111111111011",
    "1111111111110010",
    "1111111111101010",
    "1111111111100100",
    "1111111111011111",
    "1111111111011011",
    "1111111111011011",
    "1111111111011011",
    "1111111111011101",
    "1111111111011111",
    "1111111111011111",
    "1111111111011111",
    "1111111111011111",
    "1111111111011101",
    "1111111111011101",
    "1111111111011011",
    "1111111111011011",
    "1111111111011101",
    "1111111111100000",
    "1111111111100100",
    "1111111111101010",
    "1111111111101111",
    "1111111111110111",
    "1111111111111100",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111101001",
    "1111111111101010",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111111001",
    "1111111111111110",
    "0000000000000100",
    "0000000000000111",
    "0000000000000111",
    "0000000000000111",
    "0000000000000010",
    "1111111111111011",
    "1111111111110100",
    "1111111111101111",
    "1111111111101100",
    "1111111111101010",
    "1111111111101100",
    "1111111111110001",
    "1111111111111001",
    "0000000000000101",
    "0000000000010011",
    "0000000000011110",
    "0000000000101001",
    "0000000000110010",
    "0000000000110111",
    "0000000000110111",
    "0000000000110101",
    "0000000000101110",
    "0000000000100110",
    "0000000000011110",
    "0000000000010011",
    "0000000000001001",
    "1111111111111100",
    "1111111111110001",
    "1111111111100111",
    "1111111111011111",
    "1111111111011000",
    "1111111111010111",
    "1111111111011000",
    "1111111111011101",
    "1111111111100100",
    "1111111111101100",
    "1111111111110010",
    "1111111111111001",
    "0000000000000000",
    "0000000000000101",
    "0000000000001010",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010011",
    "0000000000010011",
    "0000000000010001",
    "0000000000010001",
    "0000000000010001",
    "0000000000010011",
    "0000000000010110",
    "0000000000011001",
    "0000000000011011",
    "0000000000011100",
    "0000000000011100",
    "0000000000011011",
    "0000000000010111",
    "0000000000010011",
    "0000000000001111",
    "0000000000001010",
    "0000000000000111",
    "0000000000000101",
    "0000000000000100",
    "0000000000000010",
    "0000000000000000",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101001",
    "1111111111100111",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101101",
    "1111111111110010",
    "1111111111111001",
    "0000000000000010",
    "0000000000001010",
    "0000000000010011",
    "0000000000010111",
    "0000000000011001",
    "0000000000010111",
    "0000000000010011",
    "0000000000001110",
    "0000000000000101",
    "1111111111111100",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111100",
    "0000000000000100",
    "0000000000001001",
    "0000000000001110",
    "0000000000010011",
    "0000000000010111",
    "0000000000011011",
    "0000000000011110",
    "0000000000100000",
    "0000000000100000",
    "0000000000011110",
    "0000000000011001",
    "0000000000010011",
    "0000000000001010",
    "0000000000000100",
    "1111111111111100",
    "1111111111111001",
    "1111111111111011",
    "0000000000000010",
    "0000000000001001",
    "0000000000010001",
    "0000000000011001",
    "0000000000100001",
    "0000000000101000",
    "0000000000101101",
    "0000000000101110",
    "0000000000110000",
    "0000000000110000",
    "0000000000101110",
    "0000000000101011",
    "0000000000101011",
    "0000000000101001",
    "0000000000101011",
    "0000000000101011",
    "0000000000101110",
    "0000000000110000",
    "0000000000110000",
    "0000000000110000",
    "0000000000101110",
    "0000000000101001",
    "0000000000100011",
    "0000000000011011",
    "0000000000010100",
    "0000000000001110",
    "0000000000001001",
    "0000000000000111",
    "0000000000000111",
    "0000000000001001",
    "0000000000001010",
    "0000000000001111",
    "0000000000010011",
    "0000000000010110",
    "0000000000011001",
    "0000000000011001",
    "0000000000011001",
    "0000000000010110",
    "0000000000010011",
    "0000000000001111",
    "0000000000001010",
    "0000000000000101",
    "0000000000000010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "0000000000000101",
    "0000000000001110",
    "0000000000011001",
    "0000000000100110",
    "0000000000110011",
    "0000000000111111",
    "0000000001001001",
    "0000000001001110",
    "0000000001001110",
    "0000000001001001",
    "0000000001000000",
    "0000000000110101",
    "0000000000101000",
    "0000000000011001",
    "0000000000001010",
    "1111111111111011",
    "1111111111110010",
    "1111111111101100",
    "1111111111101010",
    "1111111111101010",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000100",
    "0000000000000100",
    "0000000000000000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000001001",
    "0000000000001110",
    "0000000000010001",
    "0000000000010011",
    "0000000000010100",
    "0000000000010100",
    "0000000000010011",
    "0000000000001111",
    "0000000000001010",
    "0000000000000111",
    "0000000000000010",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111101111",
    "1111111111101010",
    "1111111111100111",
    "1111111111100100",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100101",
    "1111111111100111",
    "1111111111101100",
    "1111111111110001",
    "1111111111110110",
    "1111111111111011",
    "1111111111111110",
    "0000000000000000",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100100",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100100",
    "1111111111100111",
    "1111111111101001",
    "1111111111101100",
    "1111111111101101",
    "1111111111101101",
    "1111111111101100",
    "1111111111100111",
    "1111111111100000",
    "1111111111011010",
    "1111111111010011",
    "1111111111001110",
    "1111111111001001",
    "1111111111001001",
    "1111111111001101",
    "1111111111010000",
    "1111111111010111",
    "1111111111011111",
    "1111111111101001",
    "1111111111110010",
    "1111111111111011",
    "0000000000000101",
    "0000000000001100",
    "0000000000001111",
    "0000000000010001",
    "0000000000001111",
    "0000000000001100",
    "0000000000000111",
    "0000000000000010",
    "1111111111111011",
    "1111111111110111",
    "1111111111110010",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111100101",
    "1111111111100000",
    "1111111111011010",
    "1111111111010011",
    "1111111111001110",
    "1111111111001011",
    "1111111111001001",
    "1111111111001001",
    "1111111111001110",
    "1111111111010011",
    "1111111111011010",
    "1111111111100010",
    "1111111111101010",
    "1111111111110001",
    "1111111111110111",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111111001",
    "0000000000000101",
    "0000000000010011",
    "0000000000100011",
    "0000000000110011",
    "0000000001000100",
    "0000000001010001",
    "0000000001011100",
    "0000000001100011",
    "0000000001100110",
    "0000000001100110",
    "0000000001100001",
    "0000000001011001",
    "0000000001001110",
    "0000000000111111",
    "0000000000101110",
    "0000000000011100",
    "0000000000001100",
    "1111111111111001",
    "1111111111101001",
    "1111111111011011",
    "1111111111010000",
    "1111111111000110",
    "1111111111000001",
    "1111111110111110",
    "1111111111000001",
    "1111111111000110",
    "1111111111001101",
    "1111111111010101",
    "1111111111011010",
    "1111111111011111",
    "1111111111100010",
    "1111111111100100",
    "1111111111100100",
    "1111111111100101",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101001",
    "1111111111101001",
    "1111111111100101",
    "1111111111100010",
    "1111111111011111",
    "1111111111011011",
    "1111111111011000",
    "1111111111010101",
    "1111111111010011",
    "1111111111010010",
    "1111111111010011",
    "1111111111010111",
    "1111111111011011",
    "1111111111100000",
    "1111111111100111",
    "1111111111101101",
    "1111111111110100",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110010",
    "1111111111101101",
    "1111111111100111",
    "1111111111100010",
    "1111111111011111",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011111",
    "1111111111011111",
    "1111111111100000",
    "1111111111100000",
    "1111111111100000",
    "1111111111011111",
    "1111111111011111",
    "1111111111011101",
    "1111111111011011",
    "1111111111011011",
    "1111111111011101",
    "1111111111011111",
    "1111111111100010",
    "1111111111100101",
    "1111111111100111",
    "1111111111101010",
    "1111111111101101",
    "1111111111110001",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "0000000000000100",
    "0000000000000101",
    "0000000000000111",
    "0000000000001010",
    "0000000000001110",
    "0000000000010001",
    "0000000000010110",
    "0000000000011011",
    "0000000000100000",
    "0000000000100101",
    "0000000000101000",
    "0000000000101001",
    "0000000000101000",
    "0000000000100110",
    "0000000000100001",
    "0000000000011011",
    "0000000000010100",
    "0000000000001100",
    "0000000000000101",
    "1111111111111100",
    "1111111111110111",
    "1111111111110110",
    "1111111111110111",
    "1111111111111100",
    "0000000000000101",
    "0000000000001110",
    "0000000000010110",
    "0000000000011100",
    "0000000000100000",
    "0000000000100000",
    "0000000000011110",
    "0000000000011011",
    "0000000000010111",
    "0000000000010011",
    "0000000000001100",
    "0000000000000101",
    "1111111111111110",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110110",
    "1111111111111011",
    "0000000000000111",
    "0000000000010100",
    "0000000000100011",
    "0000000000110000",
    "0000000000111101",
    "0000000001001001",
    "0000000001001111",
    "0000000001010010",
    "0000000001010001",
    "0000000001001010",
    "0000000001000000",
    "0000000000110101",
    "0000000000101000",
    "0000000000011011",
    "0000000000001111",
    "0000000000000101",
    "1111111111111011",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111111001",
    "1111111111111110",
    "0000000000000101",
    "0000000000001010",
    "0000000000001110",
    "0000000000010011",
    "0000000000010110",
    "0000000000011011",
    "0000000000100011",
    "0000000000101011",
    "0000000000101011",
    "0000000000010110",
    "1111111111011000",
    "1111111101101110",
    "1111111011011010",
    "1111111000101011",
    "1111110101111010",
    "1111110011011101",
    "1111110001100101",
    "1111110000011000",
    "1111101111110001",
    "1111101111101001",
    "1111101111111011",
    "1111110000101000",
    "1111110001110101",
    "1111110011100101",
    "1111110101111010",
    "1111111000101011",
    "1111111011101011",
    "1111111110100101",
    "0000000001001001",
    "0000000011000010",
    "0000000100001101",
    "0000000100110001",
    "0000000101000011",
    "0000000101010111",
    "0000000101111110",
    "0000000111000011",
    "0000001000100100",
    "0000001010010101",
    "0000001100000111",
    "0000001101110000",
    "0000001111001010",
    "0000010000011001",
    "0000010001100000",
    "0000010010100100",
    "0000010011011100",
    "0000010011111010",
    "0000010011101001",
    "0000010010011011",
    "0000010000001001",
    "0000001100111100",
    "0000001001001001",
    "0000000101001011",
    "0000000001010110",
    "1111111101110100",
    "1111111010110001",
    "1111111000001101",
    "1111110110000101",
    "1111110100100000",
    "1111110011011101",
    "1111110011000110",
    "1111110011100000",
    "1111110100110000",
    "1111110110101110",
    "1111111001001111",
    "1111111100000010",
    "1111111110110001",
    "0000000001010010",
    "0000000011011010",
    "0000000101001010",
    "0000000110101010",
    "0000001000000011",
    "0000001001011000",
    "0000001010101101",
    "0000001011111010",
    "0000001100110010",
    "0000001101010000",
    "0000001101001100",
    "0000001100110010",
    "0000001100010011",
    "0000001100000001",
    "0000001100000111",
    "0000001100100111",
    "0000001101010011",
    "0000001101110111",
    "0000001101111100",
    "0000001101010110",
    "0000001100000011",
    "0000001010001011",
    "0000000111111011",
    "0000000101100100",
    "0000000011001101",
    "0000000000110111",
    "1111111110011101",
    "1111111100000000",
    "1111111001100001",
    "1111110111000111",
    "1111110101000010",
    "1111110011100010",
    "1111110010110100",
    "1111110010111100",
    "1111110011111010",
    "1111110101100000",
    "1111110111100001",
    "1111111001110000",
    "1111111100000010",
    "1111111110010010",
    "0000000000100001",
    "0000000010101000",
    "0000000100101001",
    "0000000110011010",
    "0000000111110100",
    "0000001000101100",
    "0000001001000000",
    "0000001000110001",
    "0000001000001110",
    "0000000111100101",
    "0000000111000101",
    "0000000110110100",
    "0000000110110110",
    "0000000110111101",
    "0000000111000000",
    "0000000110110001",
    "0000000110001000",
    "0000000101001010",
    "0000000011111011",
    "0000000010100110",
    "0000000001001110",
    "1111111111110010",
    "1111111110010011",
    "1111111100101001",
    "1111111010110000",
    "1111111000101011",
    "1111110110100110",
    "1111110100101101",
    "1111110011010001",
    "1111110010011101",
    "1111110010010001",
    "1111110010101010",
    "1111110011011101",
    "1111110100011011",
    "1111110101011001",
    "1111110110010110",
    "1111110111001111",
    "1111111000001100",
    "1111111001001111",
    "1111111010011100",
    "1111111011110001",
    "1111111101001000",
    "1111111110011010",
    "1111111111100000",
    "0000000000011011",
    "0000000001000100",
    "0000000001100000",
    "0000000001110010",
    "0000000001111101",
    "0000000010000100",
    "0000000010000000",
    "0000000001110101",
    "0000000001100000",
    "0000000001000000",
    "0000000000011011",
    "1111111111101101",
    "1111111110111110",
    "1111111110001101",
    "1111111101011010",
    "1111111100100111",
    "1111111011111001",
    "1111111011001111",
    "1111111010101110",
    "1111111010010101",
    "1111111010000101",
    "1111111001111110",
    "1111111001111010",
    "1111111001110110",
    "1111111001110000",
    "1111111001100110",
    "1111111001011100",
    "1111111001010110",
    "1111111001011001",
    "1111111001101011",
    "1111111010001100",
    "1111111010111011",
    "1111111011110100",
    "1111111100101110",
    "1111111101100001",
    "1111111110000110",
    "1111111110011101",
    "1111111110101001",
    "1111111110101111",
    "1111111110110111",
    "1111111111001000",
    "1111111111011111",
    "1111111111110100",
    "0000000000000101",
    "0000000000000010",
    "1111111111100111",
    "1111111110111011",
    "1111111110000011",
    "1111111101001000",
    "1111111100010100",
    "1111111011101110",
    "1111111011011100",
    "1111111011010111",
    "1111111011011100",
    "1111111011100111",
    "1111111011101110",
    "1111111011101110",
    "1111111011100010",
    "1111111011001111",
    "1111111010110110",
    "1111111010100001",
    "1111111010011001",
    "1111111010100011",
    "1111111010111110",
    "1111111011101100",
    "1111111100011111",
    "1111111101001111",
    "1111111101110110",
    "1111111110001110",
    "1111111110011101",
    "1111111110100111",
    "1111111110110100",
    "1111111111001001",
    "1111111111100101",
    "0000000000000111",
    "0000000000100011",
    "0000000000110101",
    "0000000000111010",
    "0000000000110000",
    "0000000000011001",
    "1111111111111001",
    "1111111111011011",
    "1111111111000110",
    "1111111110111100",
    "1111111111000011",
    "1111111111010011",
    "1111111111101010",
    "0000000000000100",
    "0000000000010110",
    "0000000000100000",
    "0000000000100000",
    "0000000000011001",
    "0000000000010001",
    "0000000000001001",
    "0000000000000100",
    "1111111111111110",
    "1111111111111110",
    "0000000000000010",
    "0000000000000100",
    "0000000000000111",
    "0000000000001100",
    "0000000000010001",
    "0000000000010110",
    "0000000000100000",
    "0000000000101011",
    "0000000000111000",
    "0000000001001001",
    "0000000001010110",
    "0000000001011001",
    "0000000001001111",
    "0000000000111000",
    "0000000000010001",
    "1111111111011011",
    "1111111110100010",
    "1111111101101001",
    "1111111100111000",
    "1111111100010111",
    "1111111100001011",
    "1111111100010000",
    "1111111100011111",
    "1111111100101100",
    "1111111100101110",
    "1111111100100100",
    "1111111100010100",
    "1111111100001000",
    "1111111100001000",
    "1111111100011100",
    "1111111101000001",
    "1111111101111000",
    "1111111110110111",
    "1111111111111001",
    "0000000000111000",
    "0000000001101101",
    "0000000010010100",
    "0000000010110000",
    "0000000011000000",
    "0000000011001100",
    "0000000011010111",
    "0000000011100100",
    "0000000011110101",
    "0000000100000111",
    "0000000100010101",
    "0000000100011110",
    "0000000100011001",
    "0000000100000111",
    "0000000011100110",
    "0000000010111111",
    "0000000010010100",
    "0000000001110010",
    "0000000001011110",
    "0000000001011001",
    "0000000001100011",
    "0000000001110010",
    "0000000001111010",
    "0000000001110101",
    "0000000001100000",
    "0000000000111000",
    "0000000000001100",
    "1111111111100010",
    "1111111111001000",
    "1111111111000000",
    "1111111111001001",
    "1111111111011111",
    "1111111111111001",
    "0000000000010011",
    "0000000000100110",
    "0000000000110111",
    "0000000001001010",
    "0000000001100100",
    "0000000010000111",
    "0000000010110011",
    "0000000011100110",
    "0000000100011001",
    "0000000101000111",
    "0000000101101110",
    "0000000110001101",
    "0000000110100100",
    "0000000110110110",
    "0000000111000011",
    "0000000111001101",
    "0000000111001111",
    "0000000111000101",
    "0000000110101110",
    "0000000110000011",
    "0000000101000010",
    "0000000011101001",
    "0000000001111000",
    "1111111111110010",
    "1111111101100111",
    "1111111011100100",
    "1111111001111011",
    "1111111000111101",
    "1111111000110000",
    "1111111001011001",
    "1111111010110101",
    "1111111100111000",
    "1111111111010011",
    "0000000001111010",
    "0000000100011001",
    "0000000110100010",
    "0000001000001110",
    "0000001001011010",
    "0000001010001000",
    "0000001010011010",
    "0000001010011010",
    "0000001010010000",
    "0000001010000100",
    "0000001001111100",
    "0000001001111100",
    "0000001010001001",
    "0000001010100000",
    "0000001011000001",
    "0000001011100111",
    "0000001100001110",
    "0000001100101101",
    "0000001100111110",
    "0000001100110101",
    "0000001100001011",
    "0000001010111001",
    "0000001001000001",
    "0000000110101001",
    "0000000011111110",
    "0000000001001110",
    "1111111110100010",
    "1111111100010000",
    "1111111010011100",
    "1111111001000111",
    "1111111000010001",
    "1111110111110101",
    "1111110111101001",
    "1111110111101001",
    "1111110111101000",
    "1111110111100011",
    "1111110111010110",
    "1111110111000000",
    "1111110110101001",
    "1111110110010011",
    "1111110110000101",
    "1111110110000001",
    "1111110110001100",
    "1111110110100110",
    "1111110111010001",
    "1111111000001001",
    "1111111001001111",
    "1111111010011111",
    "1111111011110001",
    "1111111101000001",
    "1111111110000101",
    "1111111110110111",
    "1111111111010011",
    "1111111111010011",
    "1111111110111001",
    "1111111110000101",
    "1111111100111101",
    "1111111011101100",
    "1111111010100001",
    "1111111001101011",
    "1111111001010110",
    "1111111001101011",
    "1111111010101011",
    "1111111100001111",
    "1111111110001010",
    "0000000000001111",
    "0000000010001100",
    "0000000011110011",
    "0000000101000000",
    "0000000101110000",
    "0000000101111110",
    "0000000101101110",
    "0000000101000010",
    "0000000011111101",
    "0000000010100100",
    "0000000001000000",
    "1111111111011010",
    "1111111101111110",
    "1111111100111000",
    "1111111100001011",
    "1111111100000000",
    "1111111100001111",
    "1111111100110100",
    "1111111101100111",
    "1111111110011101",
    "1111111111010000",
    "1111111111111011",
    "0000000000011100",
    "0000000000110011",
    "0000000001000010",
    "0000000001001110",
    "0000000001010111",
    "0000000001100000",
    "0000000001100110",
    "0000000001101110",
    "0000000001110011",
    "0000000001111000",
    "0000000001111011",
    "0000000001111101",
    "0000000010000000",
    "0000000010000101",
    "0000000010001101",
    "0000000010011011",
    "0000000010101101",
    "0000000011001000",
    "0000000011101110",
    "0000000100100001",
    "0000000101011111",
    "0000000110101010",
    "0000000111111100",
    "0000001001010000",
    "0000001010011101",
    "0000001011011101",
    "0000001100000110",
    "0000001100010101",
    "0000001100000011",
    "0000001011010000",
    "0000001001111100",
    "0000001000001110",
    "0000000110001011",
    "0000000011111110",
    "0000000001110010",
    "1111111111101101",
    "1111111101111001",
    "1111111100011101",
    "1111111011011010",
    "1111111010110001",
    "1111111010100100",
    "1111111010110000",
    "1111111011010010",
    "1111111100000110",
    "1111111101000101",
    "1111111110001010",
    "1111111111001110",
    "0000000000010110",
    "0000000001011001",
    "0000000010011001",
    "0000000011010100",
    "0000000100000101",
    "0000000100101011",
    "0000000101000101",
    "0000000101010010",
    "0000000101010101",
    "0000000101010100",
    "0000000101010111",
    "0000000101100100",
    "0000000110000000",
    "0000000110101001",
    "0000000111011010",
    "0000001000001101",
    "0000001000110111",
    "0000001001010011",
    "0000001001011101",
    "0000001001010010",
    "0000001000101111",
    "0000000111110111",
    "0000000110101010",
    "0000000101001011",
    "0000000011011010",
    "0000000001011001",
    "1111111111001011",
    "1111111100111011",
    "1111111010110001",
    "1111111000110110",
    "1111110111010010",
    "1111110110001111",
    "1111110101101101",
    "1111110101101010",
    "1111110110000100",
    "1111110110110011",
    "1111110111110010",
    "1111111000111010",
    "1111111010000111",
    "1111111011010101",
    "1111111100100100",
    "1111111101101111",
    "1111111110110110",
    "1111111111110100",
    "0000000000101101",
    "0000000001010111",
    "0000000001111010",
    "0000000010010111",
    "0000000010110001",
    "0000000011001000",
    "0000000011011110",
    "0000000011110000",
    "0000000011111101",
    "0000000100000101",
    "0000000100000101",
    "0000000011111110",
    "0000000011110011",
    "0000000011100100",
    "0000000011010101",
    "0000000011000111",
    "0000000010111000",
    "0000000010100011",
    "0000000010000010",
    "0000000001010100",
    "0000000000010110",
    "1111111111001011",
    "1111111101111011",
    "1111111100100111",
    "1111111011010111",
    "1111111010001100",
    "1111111001001100",
    "1111111000011011",
    "1111110111111011",
    "1111110111101110",
    "1111110111110011",
    "1111111000000111",
    "1111111000101000",
    "1111111001010110",
    "1111111010001101",
    "1111111011001000",
    "1111111100000010",
    "1111111100110001",
    "1111111101010000",
    "1111111101011101",
    "1111111101011000",
    "1111111101001011",
    "1111111100111011",
    "1111111100101111",
    "1111111100101111",
    "1111111100111011",
    "1111111101010000",
    "1111111101101111",
    "1111111110010010",
    "1111111110110010",
    "1111111111001011",
    "1111111111011010",
    "1111111111011011",
    "1111111111010010",
    "1111111110111001",
    "1111111110010101",
    "1111111101100100",
    "1111111100100111",
    "1111111011100010",
    "1111111010010101",
    "1111111001001100",
    "1111111000001010",
    "1111110111011100",
    "1111110111001001",
    "1111110111010010",
    "1111110111111010",
    "1111111000110110",
    "1111111001111110",
    "1111111011000111",
    "1111111100000110",
    "1111111100110110",
    "1111111101010011",
    "1111111101100100",
    "1111111101101100",
    "1111111101110110",
    "1111111110001000",
    "1111111110100010",
    "1111111111000011",
    "1111111111100111",
    "0000000000000111",
    "0000000000011110",
    "0000000000101001",
    "0000000000101110",
    "0000000000101011",
    "0000000000100101",
    "0000000000011001",
    "0000000000000111",
    "1111111111101101",
    "1111111111001110",
    "1111111110100101",
    "1111111101111011",
    "1111111101010010",
    "1111111100110001",
    "1111111100011111",
    "1111111100011100",
    "1111111100100100",
    "1111111100110110",
    "1111111101001010",
    "1111111101011101",
    "1111111101110001",
    "1111111110001000",
    "1111111110100100",
    "1111111111000000",
    "1111111111011010",
    "1111111111101001",
    "1111111111101010",
    "1111111111011111",
    "1111111111001001",
    "1111111110110110",
    "1111111110101110",
    "1111111110111011",
    "1111111111011011",
    "0000000000001111",
    "0000000001000101",
    "0000000001110101",
    "0000000010010001",
    "0000000010010111",
    "0000000010000101",
    "0000000001100000",
    "0000000000101101",
    "1111111111101010",
    "1111111110011111",
    "1111111101001000",
    "1111111011100111",
    "1111111010000000",
    "1111111000011001",
    "1111110110111010",
    "1111110101101111",
    "1111110100111100",
    "1111110100101000",
    "1111110100110101",
    "1111110101100001",
    "1111110110101000",
    "1111111000000000",
    "1111111001011100",
    "1111111010110011",
    "1111111011111001",
    "1111111100101011",
    "1111111101000110",
    "1111111101010000",
    "1111111101010011",
    "1111111101011000",
    "1111111101100101",
    "1111111101111110",
    "1111111110100010",
    "1111111111010000",
    "0000000000000101",
    "0000000000111000",
    "0000000001101000",
    "0000000010010001",
    "0000000010110110",
    "0000000011010111",
    "0000000011110110",
    "0000000100010111",
    "0000000100111000",
    "0000000101011001",
    "0000000101110100",
    "0000000110000110",
    "0000000110001101",
    "0000000110000101",
    "0000000101110000",
    "0000000101010010",
    "0000000100101110",
    "0000000100000101",
    "0000000011011001",
    "0000000010101001",
    "0000000001111010",
    "0000000001001100",
    "0000000000100011",
    "0000000000000111",
    "1111111111111100",
    "0000000000001110",
    "0000000000110011",
    "0000000001110000",
    "0000000010111000",
    "0000000100000101",
    "0000000101000111",
    "0000000101110000",
    "0000000101110011",
    "0000000101001111",
    "0000000100000000",
    "0000000010001111",
    "0000000000001100",
    "1111111110000011",
    "1111111100001011",
    "1111111010110001",
    "1111111001111010",
    "1111111001101011",
    "1111111010000010",
    "1111111010111000",
    "1111111100000101",
    "1111111101011101",
    "1111111110110110",
    "0000000000000111",
    "0000000001000100",
    "0000000001101101",
    "0000000001111111",
    "0000000001111111",
    "0000000001101110",
    "0000000001010010",
    "0000000000110010",
    "0000000000010001",
    "1111111111110100",
    "1111111111100111",
    "1111111111101010",
    "0000000000001100",
    "0000000001000111",
    "0000000010100001",
    "0000000100010111",
    "0000000110011010",
    "0000001000011100",
    "0000001010001001",
    "0000001011010000",
    "0000001011100101",
    "0000001011000011",
    "0000001001101111",
    "0000000111110110",
    "0000000101101001",
    "0000000011011010",
    "0000000001010111",
    "1111111111100111",
    "1111111110010011",
    "1111111101010111",
    "1111111100101111",
    "1111111100011010",
    "1111111100010100",
    "1111111100011000",
    "1111111100101001",
    "1111111100111110",
    "1111111101010010",
    "1111111101011000",
    "1111111101001101",
    "1111111100101100",
    "1111111011110110",
    "1111111010110110",
    "1111111001111000",
    "1111111001000101",
    "1111111000101011",
    "1111111000101101",
    "1111111001001111",
    "1111111010001111",
    "1111111011100100",
    "1111111101001000",
    "1111111110101110",
    "0000000000001100",
    "0000000001001111",
    "0000000001110110",
    "0000000001111011",
    "0000000001100011",
    "0000000000110000",
    "1111111111101100",
    "1111111110100111",
    "1111111101101100",
    "1111111101000101",
    "1111111100110100",
    "1111111100111011",
    "1111111101010011",
    "1111111101111001",
    "1111111110100111",
    "1111111111010101",
    "0000000000000101",
    "0000000000101110",
    "0000000001010100",
    "0000000001110010",
    "0000000010000100",
    "0000000010000100",
    "0000000001101110",
    "0000000001000010",
    "0000000000000100",
    "1111111110110111",
    "1111111101101010",
    "1111111100101011",
    "1111111011111110",
    "1111111011101100",
    "1111111011111000",
    "1111111100011010",
    "1111111101001111",
    "1111111110001101",
    "1111111111001101",
    "0000000000001110",
    "0000000001000111",
    "0000000001111011",
    "0000000010101110",
    "0000000011011100",
    "0000000100000101",
    "0000000100100100",
    "0000000100110011",
    "0000000100101110",
    "0000000100010010",
    "0000000011100110",
    "0000000010101001",
    "0000000001101000",
    "0000000000101011",
    "1111111111111100",
    "1111111111100111",
    "1111111111101101",
    "0000000000010011",
    "0000000001001010",
    "0000000010001111",
    "0000000011011010",
    "0000000100100010",
    "0000000101100010",
    "0000000110010101",
    "0000000110111101",
    "0000000111010101",
    "0000000111100101",
    "0000000111101111",
    "0000000111111001",
    "0000001000000000",
    "0000001000000011",
    "0000001000000011",
    "0000000111111110",
    "0000000111110100",
    "0000000111101010",
    "0000000111100010",
    "0000000111011111",
    "0000000111100001",
    "0000000111100111",
    "0000000111101110",
    "0000000111110001",
    "0000000111101100",
    "0000000111011101",
    "0000000111000011",
    "0000000110011100",
    "0000000101101110",
    "0000000100111101",
    "0000000100001100",
    "0000000011100001",
    "0000000010111000",
    "0000000010010110",
    "0000000001110011",
    "0000000001010001",
    "0000000000110000",
    "0000000000010011",
    "1111111111111001",
    "1111111111101001",
    "1111111111100101",
    "1111111111101101",
    "0000000000000111",
    "0000000000101110",
    "0000000001100110",
    "0000000010110001",
    "0000000100001010",
    "0000000101101011",
    "0000000111001010",
    "0000001000100000",
    "0000001001100111",
    "0000001010010101",
    "0000001010101101",
    "0000001010110010",
    "0000001010100111",
    "0000001010010000",
    "0000001001110001",
    "0000001001001001",
    "0000001000011000",
    "0000000111011010",
    "0000000110010000",
    "0000000100111011",
    "0000000011100011",
    "0000000010001101",
    "0000000001000100",
    "0000000000001110",
    "1111111111100111",
    "1111111111010011",
    "1111111111001101",
    "1111111111001101",
    "1111111111010000",
    "1111111111010011",
    "1111111111011000",
    "1111111111100000",
    "1111111111101111",
    "0000000000000101",
    "0000000000011110",
    "0000000000110101",
    "0000000001000111",
    "0000000001001100",
    "0000000001000100",
    "0000000000101110",
    "0000000000010011",
    "1111111111110111",
    "1111111111101001",
    "1111111111101101",
    "0000000000000111",
    "0000000000110010",
    "0000000001101001",
    "0000000010100011",
    "0000000011010111",
    "0000000011111011",
    "0000000100001010",
    "0000000100000101",
    "0000000011101100",
    "0000000011000111",
    "0000000010010110",
    "0000000001100000",
    "0000000000100000",
    "1111111111010101",
    "1111111110000011",
    "1111111100101110",
    "1111111011011001",
    "1111111010001111",
    "1111111001011001",
    "1111111000111010",
    "1111111000110011",
    "1111111001000000",
    "1111111001011010",
    "1111111001111000",
    "1111111010010010",
    "1111111010100111",
    "1111111010110011",
    "1111111010110110",
    "1111111010110110",
    "1111111010110101",
    "1111111010110101",
    "1111111010110110",
    "1111111011000000",
    "1111111011010100",
    "1111111011110100",
    "1111111100100110",
    "1111111101100101",
    "1111111110101111",
    "1111111111111011",
    "0000000001000000",
    "0000000001110101",
    "0000000010010110",
    "0000000010011110",
    "0000000010010010",
    "0000000001111000",
    "0000000001010100",
    "0000000000101110",
    "0000000000001001",
    "1111111111100010",
    "1111111111000001",
    "1111111110100010",
    "1111111110000011",
    "1111111101100001",
    "1111111100111110",
    "1111111100011000",
    "1111111011110100",
    "1111111011010100",
    "1111111010110110",
    "1111111010011001",
    "1111111001111101",
    "1111111001011110",
    "1111111000111101",
    "1111111000011100",
    "1111111000000000",
    "1111110111110000",
    "1111110111110000",
    "1111111000000010",
    "1111111000101000",
    "1111111001011100",
    "1111111010011100",
    "1111111011100001",
    "1111111100100100",
    "1111111101100100",
    "1111111110011100",
    "1111111111001011",
    "1111111111110010",
    "0000000000010110",
    "0000000000110010",
    "0000000001001001",
    "0000000001011110",
    "0000000001101110",
    "0000000001111011",
    "0000000010000100",
    "0000000010000111",
    "0000000010001000",
    "0000000010001100",
    "0000000010010001",
    "0000000010010111",
    "0000000010011100",
    "0000000010011011",
    "0000000010001000",
    "0000000001100001",
    "0000000000100011",
    "1111111111001001",
    "1111111101011111",
    "1111111011100111",
    "1111111001101110",
    "1111110111111011",
    "1111110110011011",
    "1111110101010011",
    "1111110100101000",
    "1111110100011110",
    "1111110100110000",
    "1111110101011011",
    "1111110110011001",
    "1111110111100100",
    "1111111000110110",
    "1111111010001000",
    "1111111011010100",
    "1111111100010010",
    "1111111100111101",
    "1111111101010010",
    "1111111101010000",
    "1111111100111101",
    "1111111100011101",
    "1111111011111011",
    "1111111011011111",
    "1111111011001101",
    "1111111011001011",
    "1111111011011001",
    "1111111011110100",
    "1111111100011101",
    "1111111101001111",
    "1111111110001000",
    "1111111111000110",
    "0000000000001010",
    "0000000001001010",
    "0000000010000100",
    "0000000010110001",
    "0000000011001101",
    "0000000011010100",
    "0000000011000011",
    "0000000010011011",
    "0000000001011100",
    "0000000000001001",
    "1111111110100010",
    "1111111100110110",
    "1111111011001000",
    "1111111001011111",
    "1111111000000100",
    "1111110110111111",
    "1111110110010110",
    "1111110110001100",
    "1111110110100101",
    "1111110111011100",
    "1111111000101101",
    "1111111010001101",
    "1111111011110001",
    "1111111101001101",
    "1111111110010111",
    "1111111111001000",
    "1111111111011101",
    "1111111111011011",
    "1111111111001001",
    "1111111110101100",
    "1111111110001101",
    "1111111101110011",
    "1111111101100010",
    "1111111101100001",
    "1111111101110011",
    "1111111110011010",
    "1111111111010111",
    "0000000000101011",
    "0000000010001100",
    "0000000011110011",
    "0000000101010111",
    "0000000110101110",
    "0000000111101100",
    "0000001000001110",
    "0000001000010000",
    "0000000111110011",
    "0000000110111011",
    "0000000101110000",
    "0000000100011010",
    "0000000011000010",
    "0000000001101011",
    "0000000000011110",
    "1111111111011101",
    "1111111110110010",
    "1111111110100000",
    "1111111110100101",
    "1111111111000000",
    "1111111111101010",
    "0000000000011110",
    "0000000001001111",
    "0000000001111000",
    "0000000010010100",
    "0000000010011100",
    "0000000010010001",
    "0000000001110110",
    "0000000001010010",
    "0000000000101110",
    "0000000000001110",
    "1111111111111001",
    "1111111111110110",
    "0000000000001001",
    "0000000000101011",
    "0000000001011110",
    "0000000010011011",
    "0000000011011010",
    "0000000100010101",
    "0000000101000111",
    "0000000101101011",
    "0000000101111011",
    "0000000101111011",
    "0000000101101011",
    "0000000101001101",
    "0000000100100111",
    "0000000011111101",
    "0000000011010010",
    "0000000010101101",
    "0000000010001111",
    "0000000001111000",
    "0000000001101001",
    "0000000001100000",
    "0000000001010110",
    "0000000001001001",
    "0000000000110011",
    "0000000000010011",
    "1111111111100010",
    "1111111110101100",
    "1111111101101100",
    "1111111100101110",
    "1111111011110100",
    "1111111011001000",
    "1111111010101100",
    "1111111010100011",
    "1111111010101110",
    "1111111011001010",
    "1111111011110011",
    "1111111100100100",
    "1111111101011000",
    "1111111110001010",
    "1111111110110111",
    "1111111111011011",
    "1111111111110111",
    "0000000000001100",
    "0000000000010110",
    "0000000000011011",
    "0000000000011100",
    "0000000000011011",
    "0000000000011001",
    "0000000000010110",
    "0000000000010011",
    "0000000000010001",
    "0000000000010001",
    "0000000000010110",
    "0000000000100001",
    "0000000000110111",
    "0000000001010100",
    "0000000001111010",
    "0000000010100001",
    "0000000011000111",
    "0000000011100110",
    "0000000011111010",
    "0000000100000000",
    "0000000011110110",
    "0000000011011110",
    "0000000010110110",
    "0000000010000100",
    "0000000001000111",
    "0000000000000101",
    "1111111110111110",
    "1111111101111001",
    "1111111100111011",
    "1111111100000110",
    "1111111011100010",
    "1111111011010000",
    "1111111011010101",
    "1111111011101110",
    "1111111100011000",
    "1111111101001011",
    "1111111101111110",
    "1111111110101001",
    "1111111111000101",
    "1111111111010000",
    "1111111111001101",
    "1111111110111110",
    "1111111110101001",
    "1111111110010000",
    "1111111101111001",
    "1111111101100100",
    "1111111101010011",
    "1111111101001000",
    "1111111101000101",
    "1111111101001011",
    "1111111101011111",
    "1111111101111110",
    "1111111110101100",
    "1111111111100100",
    "0000000000100011",
    "0000000001100001",
    "0000000010011100",
    "0000000011001111",
    "0000000011110110",
    "0000000100010000",
    "0000000100011001",
    "0000000100010010",
    "0000000011111101",
    "0000000011011100",
    "0000000010110001",
    "0000000010000100",
    "0000000001010110",
    "0000000000110000",
    "0000000000010111",
    "0000000000001100",
    "0000000000001111",
    "0000000000100000",
    "0000000000111101",
    "0000000001100001",
    "0000000010001000",
    "0000000010110000",
    "0000000011010100",
    "0000000011110000",
    "0000000100000011",
    "0000000100001100",
    "0000000100000101",
    "0000000011110011",
    "0000000011010100",
    "0000000010101000",
    "0000000001110000",
    "0000000000110000",
    "1111111111101100",
    "1111111110101111",
    "1111111110000000",
    "1111111101100010",
    "1111111101011111",
    "1111111101110100",
    "1111111110100000",
    "1111111111011111",
    "0000000000101011",
    "0000000001111000",
    "0000000011000011",
    "0000000100001101",
    "0000000101010100",
    "0000000110010111",
    "0000000111010011",
    "0000001000001000",
    "0000001000101100",
    "0000001000111011",
    "0000001000110010",
    "0000001000010111",
    "0000000111101001",
    "0000000110110100",
    "0000000110000011",
    "0000000101011111",
    "0000000101001010",
    "0000000101000011",
    "0000000101001000",
    "0000000101010000",
    "0000000101010111",
    "0000000101010100",
    "0000000101000101",
    "0000000100101011",
    "0000000100001000",
    "0000000011100001",
    "0000000010110110",
    "0000000010001100",
    "0000000001100001",
    "0000000000111000",
    "0000000000010001",
    "1111111111100111",
    "1111111111000001",
    "1111111110100000",
    "1111111110001000",
    "1111111101111100",
    "1111111101111100",
    "1111111110001000",
    "1111111110100000",
    "1111111111000011",
    "1111111111101101",
    "0000000000100011",
    "0000000001011110",
    "0000000010100001",
    "0000000011101001",
    "0000000100110101",
    "0000000101111110",
    "0000000110111110",
    "0000000111110001",
    "0000001000010011",
    "0000001000100010",
    "0000001000100000",
    "0000001000010000",
    "0000000111110011",
    "0000000111001011",
    "0000000110011101",
    "0000000101101001",
    "0000000100110000",
    "0000000011110000",
    "0000000010101101",
    "0000000001101001",
    "0000000000100101",
    "1111111111100010",
    "1111111110100101",
    "1111111101101100",
    "1111111100111000",
    "1111111100000101",
    "1111111011010101",
    "1111111010101001",
    "1111111010000011",
    "1111111001100100",
    "1111111001010010",
    "1111111001001111",
    "1111111001011100",
    "1111111001111010",
    "1111111010100011",
    "1111111011010101",
    "1111111100001011",
    "1111111101000101",
    "1111111110000000",
    "1111111110111100",
    "1111111111111100",
    "0000000001000000",
    "0000000010000010",
    "0000000011000000",
    "0000000011110110",
    "0000000100100001",
    "0000000100111001",
    "0000000101000010",
    "0000000100111011",
    "0000000100100111",
    "0000000100001111",
    "0000000011110011",
    "0000000011011010",
    "0000000011000101",
    "0000000010110011",
    "0000000010100011",
    "0000000010010010",
    "0000000001111101",
    "0000000001100001",
    "0000000000111101",
    "0000000000010001",
    "1111111111011101",
    "1111111110101001",
    "1111111101110100",
    "1111111101000000",
    "1111111100010000",
    "1111111011100100",
    "1111111010111110",
    "1111111010100001",
    "1111111010001101",
    "1111111010000011",
    "1111111010000011",
    "1111111010001111",
    "1111111010100100",
    "1111111010111110",
    "1111111011011111",
    "1111111100000011",
    "1111111100101011",
    "1111111101010011",
    "1111111101111100",
    "1111111110101010",
    "1111111111011011",
    "0000000000010001",
    "0000000001000111",
    "0000000001111011",
    "0000000010101101",
    "0000000011010111",
    "0000000011110011",
    "0000000100000000",
    "0000000011111010",
    "0000000011011110",
    "0000000010110001",
    "0000000001111000",
    "0000000000110011",
    "1111111111100111",
    "1111111110011101",
    "1111111101010111",
    "1111111100010101",
    "1111111011011100",
    "1111111010101110",
    "1111111010001100",
    "1111111001110101",
    "1111111001100110",
    "1111111001011110",
    "1111111001011001",
    "1111111001010111",
    "1111111001011001",
    "1111111001011110",
    "1111111001101001",
    "1111111001111101",
    "1111111010010100",
    "1111111010101110",
    "1111111011000101",
    "1111111011011001",
    "1111111011100100",
    "1111111011101001",
    "1111111011101011",
    "1111111011101100",
    "1111111011110110",
    "1111111100001010",
    "1111111100101100",
    "1111111101011010",
    "1111111110010011",
    "1111111111010011",
    "0000000000010110",
    "0000000001010001",
    "0000000010000010",
    "0000000010101001",
    "0000000011000101",
    "0000000011010101",
    "0000000011011100",
    "0000000011010111",
    "0000000011000111",
    "0000000010101101",
    "0000000010000111",
    "0000000001011011",
    "0000000000101011",
    "1111111111110111",
    "1111111111001000",
    "1111111110011111",
    "1111111101111001",
    "1111111101011000",
    "1111111100111001",
    "1111111100011010",
    "1111111011111101",
    "1111111011100001",
    "1111111011001000",
    "1111111010110011",
    "1111111010100011",
    "1111111010011001",
    "1111111010010100",
    "1111111010010100",
    "1111111010010101",
    "1111111010011010",
    "1111111010100001",
    "1111111010100111",
    "1111111010110001",
    "1111111010111110",
    "1111111011001101",
    "1111111011100001",
    "1111111011110100",
    "1111111100001000",
    "1111111100011000",
    "1111111100100001",
    "1111111100100010",
    "1111111100011101",
    "1111111100010010",
    "1111111100000000",
    "1111111011101100",
    "1111111011010101",
    "1111111010111110",
    "1111111010101001",
    "1111111010011100",
    "1111111010010101",
    "1111111010011100",
    "1111111010101011",
    "1111111011000010",
    "1111111011011111",
    "1111111100000000",
    "1111111100100100",
    "1111111101001010",
    "1111111101110100",
    "1111111110100100",
    "1111111111011011",
    "0000000000011001",
    "0000000001010010",
    "0000000010000111",
    "0000000010101110",
    "0000000011000010",
    "0000000010111111",
    "0000000010100011",
    "0000000001110011",
    "0000000000110011",
    "1111111111101001",
    "1111111110100000",
    "1111111101100001",
    "1111111100101111",
    "1111111100001111",
    "1111111100000101",
    "1111111100001101",
    "1111111100100111",
    "1111111101001101",
    "1111111101111000",
    "1111111110100111",
    "1111111111011000",
    "0000000000001110",
    "0000000001000010",
    "0000000001111010",
    "0000000010110001",
    "0000000011101001",
    "0000000100011110",
    "0000000101001010",
    "0000000101101100",
    "0000000110000011",
    "0000000110001111",
    "0000000110001101",
    "0000000101111110",
    "0000000101100110",
    "0000000101000010",
    "0000000100010101",
    "0000000011100011",
    "0000000010110000",
    "0000000010000000",
    "0000000001011001",
    "0000000000111011",
    "0000000000101011",
    "0000000000100011",
    "0000000000100001",
    "0000000000100011",
    "0000000000100101",
    "0000000000100110",
    "0000000000100110",
    "0000000000100101",
    "0000000000100110",
    "0000000000101000",
    "0000000000101001",
    "0000000000101011",
    "0000000000101011",
    "0000000000101101",
    "0000000000101101",
    "0000000000110000",
    "0000000000111010",
    "0000000001001001",
    "0000000001100000",
    "0000000001111010",
    "0000000010010111",
    "0000000010110001",
    "0000000011001000",
    "0000000011011010",
    "0000000011101000",
    "0000000011110001",
    "0000000011111101",
    "0000000100001010",
    "0000000100011010",
    "0000000100101100",
    "0000000100111101",
    "0000000101001010",
    "0000000101010000",
    "0000000101010000",
    "0000000101001011",
    "0000000101000000",
    "0000000100110101",
    "0000000100101011",
    "0000000100100100",
    "0000000100011110",
    "0000000100010111",
    "0000000100001101",
    "0000000011111110",
    "0000000011101001",
    "0000000011001101",
    "0000000010110000",
    "0000000010010001",
    "0000000001110010",
    "0000000001010111",
    "0000000000111101",
    "0000000000100101",
    "0000000000001010",
    "1111111111101101",
    "1111111111010011",
    "1111111110111011",
    "1111111110100101",
    "1111111110010111",
    "1111111110001101",
    "1111111110000110",
    "1111111110000011",
    "1111111110000011",
    "1111111110000101",
    "1111111110001010",
    "1111111110010011",
    "1111111110100010",
    "1111111110110111",
    "1111111111010011",
    "1111111111110010",
    "0000000000010111",
    "0000000000110111",
    "0000000001010100",
    "0000000001101011",
    "0000000001111010",
    "0000000010000100",
    "0000000010000111",
    "0000000010001000",
    "0000000010001010",
    "0000000010001010",
    "0000000010001010",
    "0000000010001000",
    "0000000010000101",
    "0000000010000000",
    "0000000001111010",
    "0000000001110101",
    "0000000001110101",
    "0000000001111101",
    "0000000010001100",
    "0000000010100011",
    "0000000010111111",
    "0000000011010111",
    "0000000011101011",
    "0000000011110110",
    "0000000011110101",
    "0000000011100110",
    "0000000011001010",
    "0000000010100011",
    "0000000001110000",
    "0000000000110011",
    "1111111111101101",
    "1111111110100111",
    "1111111101100001",
    "1111111100011111",
    "1111111011100111",
    "1111111011000000",
    "1111111010110000",
    "1111111010111001",
    "1111111011011100",
    "1111111100011000",
    "1111111101100101",
    "1111111110111110",
    "0000000000010110",
    "0000000001100100",
    "0000000010100100",
    "0000000011010010",
    "0000000011110001",
    "0000000100000000",
    "0000000011111110",
    "0000000011110000",
    "0000000011010100",
    "0000000010101101",
    "0000000001111011",
    "0000000001001001",
    "0000000000010111",
    "1111111111101100",
    "1111111111001110",
    "1111111110111100",
    "1111111110110110",
    "1111111110110111",
    "1111111111000000",
    "1111111111001001",
    "1111111111010010",
    "1111111111010101",
    "1111111111010101",
    "1111111111001110",
    "1111111110111110",
    "1111111110100111",
    "1111111110001000",
    "1111111101100100",
    "1111111100111110",
    "1111111100011010",
    "1111111011111011",
    "1111111011100001",
    "1111111011001101",
    "1111111011000000",
    "1111111010111101",
    "1111111011000011",
    "1111111011010100",
    "1111111011110000",
    "1111111100011000",
    "1111111101001011",
    "1111111110001000",
    "1111111111001011",
    "0000000000010111",
    "0000000001100000",
    "0000000010101000",
    "0000000011100100",
    "0000000100010111",
    "0000000100111001",
    "0000000101001111",
    "0000000101011001",
    "0000000101011100",
    "0000000101011101",
    "0000000101011111",
    "0000000101100111",
    "0000000101110011",
    "0000000110000010",
    "0000000110010010",
    "0000000110100010",
    "0000000110110001",
    "0000000110111101",
    "0000000111000101",
    "0000000111001011",
    "0000000111001101",
    "0000000111001010",
    "0000000110111110",
    "0000000110100111",
    "0000000110000010",
    "0000000101001010",
    "0000000100000010",
    "0000000010101011",
    "0000000001001010",
    "1111111111100100",
    "1111111110000001",
    "1111111100100110",
    "1111111011010111",
    "1111111010011001",
    "1111111001101100",
    "1111111001011001",
    "1111111001011010",
    "1111111001110011",
    "1111111010100001",
    "1111111011011111",
    "1111111100101011",
    "1111111101111100",
    "1111111111010011",
    "0000000000101001",
    "0000000001110101",
    "0000000010110110",
    "0000000011101000",
    "0000000100001000",
    "0000000100010101",
    "0000000100001111",
    "0000000011111000",
    "0000000011010100",
    "0000000010101001",
    "0000000001111011",
    "0000000001010001",
    "0000000000101011",
    "0000000000001100",
    "1111111111101111",
    "1111111111011000",
    "1111111111000101",
    "1111111110110100",
    "1111111110100100",
    "1111111110010010",
    "1111111101111110",
    "1111111101100101",
    "1111111101001010",
    "1111111100100110",
    "1111111011111011",
    "1111111011000101",
    "1111111010001010",
    "1111111001000101",
    "1111110111111111",
    "1111110110111100",
    "1111110110000010",
    "1111110101011000",
    "1111110101000100",
    "1111110101001100",
    "1111110101110011",
    "1111110110110101",
    "1111111000001111",
    "1111111001111010",
    "1111111011101100",
    "1111111101011100",
    "1111111111000011",
    "0000000000011100",
    "0000000001100001",
    "0000000010010010",
    "0000000010110011",
    "0000000011000010",
    "0000000011000000",
    "0000000010110000",
    "0000000010010010",
    "0000000001101011",
    "0000000001000000",
    "0000000000011001",
    "1111111111110111",
    "1111111111100111",
    "1111111111100010",
    "1111111111100101",
    "1111111111101100",
    "1111111111101101",
    "1111111111101001",
    "1111111111011011",
    "1111111111000011",
    "1111111110100101",
    "1111111110000110",
    "1111111101100111",
    "1111111101001010",
    "1111111100110001",
    "1111111100011101",
    "1111111100001101",
    "1111111100000010",
    "1111111011111001",
    "1111111011110110",
    "1111111011111001",
    "1111111100000010",
    "1111111100010101",
    "1111111100110001",
    "1111111101011000",
    "1111111110000110",
    "1111111110111100",
    "1111111111110110",
    "0000000000110011",
    "0000000001101101",
    "0000000010100001",
    "0000000011010001",
    "0000000011110101",
    "0000000100001101",
    "0000000100010101",
    "0000000100001111",
    "0000000011111000",
    "0000000011010111",
    "0000000010101110",
    "0000000010000010",
    "0000000001010100",
    "0000000000100110",
    "1111111111110110",
    "1111111111001000",
    "1111111110011000",
    "1111111101101001",
    "1111111100111011",
    "1111111100010000",
    "1111111011101110",
    "1111111011010100",
    "1111111011000010",
    "1111111010111000",
    "1111111010110011",
    "1111111010101100",
    "1111111010100100",
    "1111111010011100",
    "1111111010010101",
    "1111111010010010",
    "1111111010010100",
    "1111111010011110",
    "1111111010101100",
    "1111111011000000",
    "1111111011010111",
    "1111111011110011",
    "1111111100010010",
    "1111111100111000",
    "1111111101100100",
    "1111111110010101",
    "1111111111001001",
    "1111111111111110",
    "0000000000110000",
    "0000000001011001",
    "0000000001111000",
    "0000000010001111",
    "0000000010011011",
    "0000000010011001",
    "0000000010001100",
    "0000000001110101",
    "0000000001010010",
    "0000000000101001",
    "1111111111111001",
    "1111111111000101",
    "1111111110001110",
    "1111111101010111",
    "1111111100011111",
    "1111111011101011",
    "1111111010111011",
    "1111111010010101",
    "1111111001111101",
    "1111111001110101",
    "1111111001111101",
    "1111111010010101",
    "1111111010111011",
    "1111111011101110",
    "1111111100100110",
    "1111111101011101",
    "1111111110010000",
    "1111111110111011",
    "1111111111011101",
    "1111111111111001",
    "0000000000010111",
    "0000000000110011",
    "0000000001010001",
    "0000000001110011",
    "0000000010010110",
    "0000000010111010",
    "0000000011011111",
    "0000000100001010",
    "0000000100111001",
    "0000000101101110",
    "0000000110100111",
    "0000000111100001",
    "0000001000010111",
    "0000001001000001",
    "0000001001011101",
    "0000001001100111",
    "0000001001100000",
    "0000001001001001",
    "0000001000100101",
    "0000000111110111",
    "0000000110111110",
    "0000000101111101",
    "0000000100110101",
    "0000000011101001",
    "0000000010011111",
    "0000000001100000",
    "0000000000101110",
    "0000000000010001",
    "0000000000001010",
    "0000000000010110",
    "0000000000110010",
    "0000000001011001",
    "0000000010000100",
    "0000000010110011",
    "0000000011100011",
    "0000000100010010",
    "0000000101000010",
    "0000000101101100",
    "0000000110010000",
    "0000000110101010",
    "0000000110111001",
    "0000000110111011",
    "0000000110110001",
    "0000000110011111",
    "0000000110001000",
    "0000000101110000",
    "0000000101011001",
    "0000000101000011",
    "0000000100110001",
    "0000000100011110",
    "0000000100001000",
    "0000000011110001",
    "0000000011010101",
    "0000000010111000",
    "0000000010011001",
    "0000000001111000",
    "0000000001010111",
    "0000000000110101",
    "0000000000010100",
    "1111111111110001",
    "1111111111010011",
    "1111111110110111",
    "1111111110100000",
    "1111111110001101",
    "1111111110000000",
    "1111111101111000",
    "1111111101110110",
    "1111111101111011",
    "1111111110000101",
    "1111111110010011",
    "1111111110100101",
    "1111111110111011",
    "1111111111001110",
    "1111111111100000",
    "1111111111110001",
    "1111111111111100",
    "0000000000000101",
    "0000000000000101",
    "1111111111111100",
    "1111111111110001",
    "1111111111100000",
    "1111111111001101",
    "1111111110111001",
    "1111111110101001",
    "1111111110011101",
    "1111111110011000",
    "1111111110011010",
    "1111111110100000",
    "1111111110101010",
    "1111111110110111",
    "1111111111001001",
    "1111111111100000",
    "1111111111111110",
    "0000000000101001",
    "0000000001011100",
    "0000000010011011",
    "0000000011011111",
    "0000000100100110",
    "0000000101101011",
    "0000000110100010",
    "0000000111001011",
    "0000000111100100",
    "0000000111101110",
    "0000000111101100",
    "0000000111100101",
    "0000000111011101",
    "0000000111010111",
    "0000000111010101",
    "0000000111010011",
    "0000000111010010",
    "0000000111001101",
    "0000000111000001",
    "0000000110101100",
    "0000000110001111",
    "0000000101100110",
    "0000000100110101",
    "0000000011110110",
    "0000000010110000",
    "0000000001100000",
    "0000000000001001",
    "1111111110101010",
    "1111111101001011",
    "1111111011101011",
    "1111111010001101",
    "1111111000110101",
    "1111110111101000",
    "1111110110101000",
    "1111110101111010",
    "1111110101100011",
    "1111110101100101",
    "1111110101111101",
    "1111110110101011",
    "1111110111101110",
    "1111111001000000",
    "1111111010011001",
    "1111111011110000",
    "1111111100111101",
    "1111111101111001",
    "1111111110011111",
    "1111111110101110",
    "1111111110100101",
    "1111111110001010",
    "1111111101100010",
    "1111111100101111",
    "1111111011111001",
    "1111111010111110",
    "1111111010000011",
    "1111111001000111",
    "1111111000001101",
    "1111110111011100",
    "1111110110110101",
    "1111110110011001",
    "1111110110001100",
    "1111110110000111",
    "1111110110001010",
    "1111110110010001",
    "1111110110011011",
    "1111110110100011",
    "1111110110101001",
    "1111110110110010",
    "1111110110110111",
    "1111110110111000",
    "1111110110110000",
    "1111110110100000",
    "1111110110000101",
    "1111110101100011",
    "1111110101000010",
    "1111110100100110",
    "1111110100011011",
    "1111110100100001",
    "1111110100111111",
    "1111110101110011",
    "1111110110111100",
    "1111111000010100",
    "1111111001111000",
    "1111111011100010",
    "1111111101001101",
    "1111111110110010",
    "0000000000010100",
    "0000000001101001",
    "0000000010110011",
    "0000000011101100",
    "0000000100010111",
    "0000000100110011",
    "0000000101000111",
    "0000000101010010",
    "0000000101011111",
    "0000000101101011",
    "0000000101110110",
    "0000000110000010",
    "0000000110001000",
    "0000000110000010",
    "0000000101101110",
    "0000000101001010",
    "0000000100010101",
    "0000000011010010",
    "0000000010001010",
    "0000000001000010",
    "1111111111111110",
    "1111111111001001",
    "1111111110100100",
    "1111111110001110",
    "1111111110000011",
    "1111111110000000",
    "1111111110000001",
    "1111111110000011",
    "1111111110000001",
    "1111111101111000",
    "1111111101100101",
    "1111111101001000",
    "1111111100011111",
    "1111111011110000",
    "1111111011000000",
    "1111111010011010",
    "1111111010000101",
    "1111111010001100",
    "1111111010110000",
    "1111111011110000",
    "1111111101000110",
    "1111111110101100",
    "0000000000011001",
    "0000000010000101",
    "0000000011101001",
    "0000000101000101",
    "0000000110010010",
    "0000000111001111",
    "0000000111111001",
    "0000001000010011",
    "0000001000011100",
    "0000001000010101",
    "0000001000000000",
    "0000000111011111",
    "0000000110110100",
    "0000000110000010",
    "0000000101001101",
    "0000000100010101",
    "0000000011100001",
    "0000000010110000",
    "0000000010000111",
    "0000000001100110",
    "0000000001001110",
    "0000000000111000",
    "0000000000100101",
    "0000000000001010",
    "1111111111100101",
    "1111111110111011",
    "1111111110001010",
    "1111111101010111",
    "1111111100100110",
    "1111111011111011",
    "1111111011011010",
    "1111111011000010",
    "1111111010110001",
    "1111111010101001",
    "1111111010100111",
    "1111111010110000",
    "1111111011000101",
    "1111111011101011",
    "1111111100100001",
    "1111111101100101",
    "1111111110110110",
    "0000000000010011",
    "0000000001101110",
    "0000000011001100",
    "0000000100100110",
    "0000000101110110",
    "0000000110110011",
    "0000000111011000",
    "0000000111100010",
    "0000000111001111",
    "0000000110100100",
    "0000000101101011",
    "0000000100110000",
    "0000000100000011",
    "0000000011110000",
    "0000000011111101",
    "0000000100101001",
    "0000000101110000",
    "0000000111001000",
    "0000001000100010",
    "0000001001110111",
    "0000001010111100",
    "0000001011101101",
    "0000001100001011",
    "0000001100010001",
    "0000001100000011",
    "0000001011100000",
    "0000001010101000",
    "0000001001100000",
    "0000001000001010",
    "0000000110101110",
    "0000000101010010",
    "0000000100000011",
