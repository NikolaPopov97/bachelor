----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/16/2022 03:00:20 PM
-- Design Name: 
-- Module Name: coef_rom - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity coef_rom is
    Port ( addr : in STD_LOGIC_VECTOR (15 downto 0);
           clk : in STD_LOGIC;
           data : out STD_LOGIC_VECTOR (15 downto 0));
end coef_rom;

architecture Behavioral of coef_rom is
type rom_type is array (22049 downto 0) of std_logic_vector(15 downto 0);

signal ROM : rom_type := 
("1100000111001101",
"1100000111001101",
"1100000111001101",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111001111",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010000",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010010",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010011",
"1100000111010101",
"1100000111010101",
"1100000111010101",
"1100000111010101",
"1100000111010101",
"1100000111010101",
"1100000111010101",
"1100000111010101",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111010111",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011000",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011010",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011100",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011101",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111011111",
"1100000111100001",
"1100000111100001",
"1100000111100001",
"1100000111100001",
"1100000111100001",
"1100000111100001",
"1100000111100001",
"1100000111100001",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100010",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100100",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100101",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111100111",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101001",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101010",
"1100000111101100",
"1100000111101100",
"1100000111101100",
"1100000111101100",
"1100000111101100",
"1100000111101100",
"1100000111101100",
"1100000111101100",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101110",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111101111",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110001",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110011",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110100",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110110",
"1100000111110111",
"1100000111110111",
"1100000111110111",
"1100000111110111",
"1100000111110111",
"1100000111110111",
"1100000111110111",
"1100000111110111",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111001",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111011",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111100",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100000111111110",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000000",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000001",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000011",
"1100001000000101",
"1100001000000101",
"1100001000000101",
"1100001000000101",
"1100001000000101",
"1100001000000101",
"1100001000000101",
"1100001000000101",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000000110",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001000",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001010",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001011",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001101",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000001110",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010000",
"1100001000010010",
"1100001000010010",
"1100001000010010",
"1100001000010010",
"1100001000010010",
"1100001000010010",
"1100001000010010",
"1100001000010010",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010011",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010101",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000010111",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011000",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011010",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011100",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011101",
"1100001000011111",
"1100001000011111",
"1100001000011111",
"1100001000011111",
"1100001000011111",
"1100001000011111",
"1100001000011111",
"1100001000011111",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100000",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100010",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100100",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100101",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000100111",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101001",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101010",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101100",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101110",
"1100001000101111",
"1100001000101111",
"1100001000101111",
"1100001000101111",
"1100001000101111",
"1100001000101111",
"1100001000101111",
"1100001000101111",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110001",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110010",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110100",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110110",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000110111",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111001",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111011",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111100",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001000111110",
"1100001001000000",
"1100001001000000",
"1100001001000000",
"1100001001000000",
"1100001001000000",
"1100001001000000",
"1100001001000000",
"1100001001000000",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000001",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000011",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000100",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001000110",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001000",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001001",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001011",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001101",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001001110",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010000",
"1100001001010010",
"1100001001010010",
"1100001001010010",
"1100001001010010",
"1100001001010010",
"1100001001010010",
"1100001001010010",
"1100001001010010",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010011",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010101",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001010111",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011000",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011010",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011011",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011101",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001011111",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100000",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100010",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100100",
"1100001001100101",
"1100001001100101",
"1100001001100101",
"1100001001100101",
"1100001001100101",
"1100001001100101",
"1100001001100101",
"1100001001100101",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001100111",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101001",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101010",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101100",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101101",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001101111",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110001",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110010",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110100",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110110",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001110111",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111001",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111011",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111100",
"1100001001111110",
"1100001001111110",
"1100001001111110",
"1100001001111110",
"1100001001111110",
"1100001001111110",
"1100001001111110",
"1100001001111110",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001001111111",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000001",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000011",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000100",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010000110",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001000",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001001",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001011",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001101",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010001110",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010000",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010001",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010011",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010101",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010010110",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011000",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011010",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011011",
"1100001010011101",
"1100001010011101",
"1100001010011101",
"1100001010011101",
"1100001010011101",
"1100001010011101",
"1100001010011101",
"1100001010011101",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010011111",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100000",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100010",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100100",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100101",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010100111",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101000",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101010",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101100",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101101",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010101111",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110001",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110010",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110100",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110110",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010110111",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111001",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111010",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111100",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111110",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001010111111",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000001",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000011",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000100",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011000110",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001000",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001001",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001011",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001100",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011001110",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010000",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010001",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010011",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010101",
"1100001011010110",
"1100001011010110",
"1100001011010110",
"1100001011010110",
"1100001011010110",
"1100001011010110",
"1100001011010110",
"1100001011010110",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011000",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011010",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011011",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011101",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011011111",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100000",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100010",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100011",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100101",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011100111",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101000",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101010",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101100",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101101",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011101111",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110001",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110010",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110100",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110101",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011110111",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111001",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111010",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111100",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111110",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001011111111",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000001",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000011",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000100",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000110",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100000111",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001001",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001011",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001100",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100001110",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010000",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010001",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010011",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010101",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100010110",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011000",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011001",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011011",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011101",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100011110",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100000",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100010",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100011",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100101",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100100111",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101000",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101010",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101100",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101101",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100101111",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110000",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110010",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110100",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110101",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100110111",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111001",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111010",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111100",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111110",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001100111111",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000001",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000010",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000100",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000110",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101000111",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001001",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001011",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001100",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101001110",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010000",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010001",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010011",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010100",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101010110",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011000",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011001",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011011",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011101",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101011110",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100000",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100010",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100011",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100101",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101100110",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101000",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101010",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101011",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101101",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101101111",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110000",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110010",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110100",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110101",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101110111",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111001",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111010",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111100",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111101",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001101111111",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000001",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000010",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000100",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000110",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110000111",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001001",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001011",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001100",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001110",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110001111",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010001",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010011",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010100",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110010110",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011000",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011001",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011011",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011101",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110011110",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100000",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100001",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100011",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100101",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110100110",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101000",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101010",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101011",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101101",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110101111",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110000",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110010",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110011",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110101",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110110111",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111000",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111010",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111100",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111101",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001110111111",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000001",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000010",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000100",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000110",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111000111",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001001",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001010",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001100",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001110",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111001111",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010001",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010011",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010100",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111010110",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011000",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011001",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011011",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011100",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111011110",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100000",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100001",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100011",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100101",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111100110",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101000",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101010",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101011",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101101",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111101110",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110000",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110010",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110011",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110101",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111110111",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111000",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111010",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111100",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111101",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100001111111111",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000001",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000010",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000100",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000101",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000000111",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001001",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001010",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001100",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001110",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000001111",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010001",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010011",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010100",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010110",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000010111",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011001",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011011",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011100",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000011110",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100000",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100001",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100011",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100101",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000100110",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101000",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101001",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101011",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101101",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000101110",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110000",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110010",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110011",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110101",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000110111",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111000",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111010",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111011",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111101",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010000111111",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000000",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000010",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000100",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000101",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001000111",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001001",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001010",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001100",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001110",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001001111",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010001",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010010",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010100",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010110",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001010111",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011001",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011011",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011100",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001011110",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100000",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100001",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100011",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100100",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001100110",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101000",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101001",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101011",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101101",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001101110",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110000",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110010",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110011",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110101",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001110110",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111000",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111010",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111011",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111101",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010001111111",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000000",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000010",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000100",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000101",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010000111",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001000",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001010",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001100",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001101",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010001111",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010001",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010010",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010100",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010110",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010010111",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011001",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011011",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011100",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011110",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010011111",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100001",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100011",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100100",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010100110",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101000",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101001",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101011",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101101",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010101110",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110000",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110001",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110011",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110101",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010110110",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111000",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111010",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111011",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111101",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010010111111",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000000",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000010",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000011",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000101",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011000111",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001000",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001010",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001100",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001101",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011001111",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010001",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010010",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010100",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010101",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011010111",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011001",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011010",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011100",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011110",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011011111",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100001",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100011",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100100",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011100110",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101000",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101001",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101011",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101100",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011101110",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110000",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110001",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110011",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110101",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011110110",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111000",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111010",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111011",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111101",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010011111110",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000000",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000010",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000011",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000101",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100000111",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001000",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001010",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001100",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001101",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100001111",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010000",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010010",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010100",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010101",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100010111",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011001",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011010",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011100",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011110",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100011111",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100001",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100010",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100100",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100110",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100100111",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101001",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101011",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101100",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100101110",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110000",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110001",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110011",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110101",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100110110",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111000",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111001",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111011",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111101",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010100111110",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000000",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000010",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000011",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000101",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101000111",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001000",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001010",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001011",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001101",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101001111",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010000",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010010",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010100",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010101",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101010111",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011001",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011010",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011100",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011101",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101011111",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100001",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100010",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100100",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100110",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101100111",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101001",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101011",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101100",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101101110",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110000",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110001",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110011",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110100",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101110110",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111000",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111001",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111011",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111101",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010101111110",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000000",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000010",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000011",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000101",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110000110",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001000",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001010",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001011",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001101",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110001111",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010000",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010010",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010100",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010101",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110010111",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011000",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011010",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011100",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011101",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110011111",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100001",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100010",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100100",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100110",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110100111",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101001",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101010",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101100",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101110",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110101111",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110001",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110011",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110100",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110110110",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111000",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111001",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111011",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111101",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010110111110",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000000",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000001",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000011",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000101",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111000110",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001000",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001010",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001011",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001101",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111001111",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010000",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010010",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010011",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010101",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111010111",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011000",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011010",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011100",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011101",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111011111",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100001",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100010",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100100",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100101",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111100111",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101001",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101010",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101100",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101110",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111101111",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110001",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110011",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110100",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110110",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111110111",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111001",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111011",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111100",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100010111111110",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000000",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000001",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000011",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000101",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000000110",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001000",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001010",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001011",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001101",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000001110",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010000",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010010",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010011",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010101",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000010111",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011000",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011010",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011100",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011101",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000011111",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100000",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100010",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100100",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100101",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000100111",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101001",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101010",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101100",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101110",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000101111",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110001",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110010",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110100",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110110",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000110111",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111001",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111011",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111100",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011000111110",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000000",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000001",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000011",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000100",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001000110",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001000",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001001",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001011",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001101",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001001110",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010000",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010010",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010011",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010101",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001010111",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011000",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011010",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011011",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011101",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001011111",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100000",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100010",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100100",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100101",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001100111",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101001",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101010",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101100",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101101",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001101111",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110001",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110010",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110100",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110110",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001110111",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111001",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111011",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111100",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111110",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011001111111",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000001",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000011",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000100",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010000110",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001000",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001001",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001011",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001101",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010001110",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010000",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010001",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010011",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010101",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010010110",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011000",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011010",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011011",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011101",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010011111",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100000",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100010",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100100",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100101",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010100111",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101000",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101010",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101100",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101101",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010101111",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110001",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110010",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110100",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110110",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010110111",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111001",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111010",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111100",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111110",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011010111111",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000001",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000011",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000100",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011000110",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001000",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001001",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001011",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001100",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011001110",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010000",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010001",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010011",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010101",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011010110",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011000",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011010",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011011",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011101",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011011111",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100000",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100010",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100011",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100101",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011100111",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101000",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101010",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101100",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101101",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011101111",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110001",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110010",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110100",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110101",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011110111",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111001",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111010",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111100",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111110",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011011111111",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000001",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000011",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000100",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000110",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100000111",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001001",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001011",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001100",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100001110",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010000",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010001",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010011",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010101",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100010110",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011000",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011001",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011011",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011101",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100011110",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100000",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100010",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100011",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100101",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100100111",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101000",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101010",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101100",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101101",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100101111",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110000",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110010",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110100",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110101",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100110111",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111001",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111010",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111100",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111110",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011100111111",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000001",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000010",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000100",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000110",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101000111",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001001",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001011",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001100",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101001110",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010000",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010001",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010011",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010100",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101010110",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011000",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011001",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011011",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011101",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101011110",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100000",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100010",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100011",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100101",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101100110",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101000",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101010",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101011",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101101",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101101111",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110000",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110010",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110100",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110101",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101110111",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111001",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111010",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111100",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111101",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011101111111",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000001",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000010",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000100",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000110",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110000111",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001001",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001011",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001100",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001110",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110001111",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010001",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010011",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010100",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110010110",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011000",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011001",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011011",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011101",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110011110",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100000",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100001",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100011",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100101",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110100110",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101000",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101010",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101011",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101101",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110101111",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110000",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110010",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110011",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110101",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110110111",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111000",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111010",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111100",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111101",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011110111111",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000001",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000010",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000100",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000110",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111000111",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001001",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001010",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001100",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001110",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111001111",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010001",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010011",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010100",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111010110",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011000",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011001",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011011",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011100",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111011110",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100000",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100001",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100011",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100101",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111100110",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101000",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101010",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101011",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101101",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111101110",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110000",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110010",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110011",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110101",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111110111",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111000",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111010",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111100",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111101",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100011111111111",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000001",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000010",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000100",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000101",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000000111",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001001",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001010",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001100",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001110",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000001111",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010001",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010011",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010100",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010110",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000010111",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011001",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011011",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011100",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000011110",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100000",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100001",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100011",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100101",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000100110",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101000",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101001",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101011",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101101",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000101110",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110000",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110010",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110011",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110101",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000110111",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111000",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111010",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111011",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111101",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100000111111",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000000",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000010",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000100",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000101",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001000111",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001001",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001010",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001100",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001110",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001001111",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010001",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010010",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010100",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010110",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001010111",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011001",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011011",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011100",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001011110",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100000",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100001",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100011",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100100",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001100110",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101000",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101001",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101011",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101101",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001101110",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110000",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110010",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110011",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110101",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001110110",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111000",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111010",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111011",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111101",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100001111111",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000000",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000010",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000100",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000101",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010000111",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001000",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001010",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001100",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001101",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010001111",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010001",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010010",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010100",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010110",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010010111",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011001",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011011",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011100",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011110",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010011111",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100001",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100011",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100100",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010100110",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101000",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101001",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101011",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101101",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010101110",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110000",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110001",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110011",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110101",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010110110",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111000",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111010",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111011",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111101",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100010111111",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000000",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000010",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000011",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000101",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011000111",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001000",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001010",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001100",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001101",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011001111",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010001",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010010",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010100",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010101",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011010111",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011001",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011010",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011100",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011110",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011011111",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100001",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100011",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100100",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011100110",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101000",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101001",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101011",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101100",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011101110",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110000",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110001",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110011",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110101",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011110110",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111000",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111010",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111011",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111101",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100011111110",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000000",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000010",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000011",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000101",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100000111",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001000",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001010",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001100",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001101",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100001111",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010000",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010010",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010100",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010101",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100010111",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011001",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011010",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011100",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011110",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100011111",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100001",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100010",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100100",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100110",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100100111",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101001",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101011",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101100",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100101110",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110000",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110001",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110011",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110101",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100110110",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111000",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111001",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111011",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111101",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100100111110",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000000",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000010",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000011",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000101",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101000111",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001000",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001010",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001011",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001101",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101001111",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010000",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010010",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010100",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010101",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101010111",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011001",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011010",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011100",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011101",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101011111",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100001",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100010",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100100",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100110",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101100111",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101001",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101011",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101100",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101101110",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110000",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110001",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110011",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110100",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101110110",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111000",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111001",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111011",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111101",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100101111110",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000000",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000010",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000011",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000101",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110000110",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001000",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001010",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001011",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001101",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110001111",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010000",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010010",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010100",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010101",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110010111",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011000",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011010",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011100",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011101",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110011111",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100001",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100010",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100100",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100110",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110100111",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101001",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101010",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101100",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101110",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110101111",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110001",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110011",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110100",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110110110",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111000",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111001",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111011",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111101",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100110111110",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000000",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000001",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000011",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000101",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111000110",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001000",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001010",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001011",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001101",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111001111",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010000",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010010",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010011",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010101",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111010111",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011000",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011010",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011100",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011101",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111011111",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100001",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100010",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100100",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100101",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111100111",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101001",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101010",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101100",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101110",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111101111",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110001",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110011",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110100",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110110",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111110111",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111001",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111011",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111100",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100100111111110",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000000",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000001",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000011",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000101",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000000110",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001000",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001010",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001011",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001101",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000001110",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010000",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010010",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010011",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010101",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000010111",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011000",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011010",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011100",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011101",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000011111",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100000",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100010",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100100",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100101",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000100111",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101001",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101010",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101100",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101110",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000101111",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110001",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110010",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110100",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110110",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000110111",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111001",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111011",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111100",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101000111110",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000000",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000001",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000011",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000100",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001000110",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001000",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001001",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001011",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001101",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001001110",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010000",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010010",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010011",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010101",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001010111",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011000",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011010",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011011",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011101",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001011111",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100000",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100010",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100100",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100101",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001100111",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101001",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101010",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101100",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101101",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001101111",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110001",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110010",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110100",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110110",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001110111",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111001",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111011",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111100",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111110",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101001111111",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000001",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000011",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000100",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010000110",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001000",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001001",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001011",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001101",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010001110",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010000",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010001",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010011",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010101",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010010110",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011000",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011010",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011011",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011101",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010011111",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100000",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100010",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100100",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100101",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010100111",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101000",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101010",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101100",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101101",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010101111",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110001",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110010",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110100",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110110",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010110111",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111001",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111010",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111100",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111110",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101010111111",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000001",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000011",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000100",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011000110",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001000",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001001",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001011",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001100",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011001110",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010000",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010001",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010011",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010101",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011010110",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011000",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011010",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011011",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011101",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011011111",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100000",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100010",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100011",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100101",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011100111",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101000",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101010",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101100",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101101",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011101111",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110001",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110010",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110100",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110101",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011110111",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111001",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111010",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111100",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111110",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101011111111",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000001",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000011",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000100",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000110",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100000111",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001001",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001011",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001100",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100001110",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010000",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010001",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010011",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010101",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100010110",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011000",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011001",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011011",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011101",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100011110",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100000",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100010",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100011",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100101",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100100111",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101000",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101010",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101100",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101101",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100101111",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110000",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110010",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110100",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110101",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100110111",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111001",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111010",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111100",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111110",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101100111111",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000001",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000010",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000100",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000110",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101000111",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001001",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001011",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001100",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101001110",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010000",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010001",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010011",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010100",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101010110",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011000",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011001",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011011",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011101",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101011110",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100000",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100010",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100011",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100101",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101100110",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101000",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101010",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101011",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101101",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101101111",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110000",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110010",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110100",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110101",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101110111",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111001",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111010",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111100",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111101",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101101111111",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000001",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000010",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000100",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000110",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110000111",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001001",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001011",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001100",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001110",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110001111",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010001",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010011",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010100",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110010110",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011000",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011001",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011011",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011101",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110011110",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100000",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100001",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100011",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100101",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110100110",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101000",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101010",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101011",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101101",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110101111",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110000",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110010",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110011",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110101",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110110111",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111000",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111010",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111100",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111101",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101110111111",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000001",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000010",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000100",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000110",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111000111",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001001",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001010",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001100",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001110",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111001111",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010001",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010011",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010100",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111010110",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011000",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011001",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011011",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011100",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111011110",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100000",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100001",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100011",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100101",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111100110",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101000",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101010",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101011",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101101",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111101110",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110000",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110010",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110011",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110101",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111110111",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111000",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111010",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111100",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111101",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100101111111111",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000001",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000010",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000100",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000101",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000000111",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001001",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001010",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001100",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001110",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000001111",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010001",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010011",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010100",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010110",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000010111",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011001",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011011",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011100",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000011110",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100000",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100001",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100011",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100101",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000100110",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101000",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101001",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101011",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101101",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000101110",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110000",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110010",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110011",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110101",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000110111",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111000",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111010",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111011",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111101",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110000111111",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000000",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000010",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000100",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000101",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001000111",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001001",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001010",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001100",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001110",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001001111",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010001",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010010",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010100",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010110",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001010111",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011001",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011011",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011100",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001011110",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100000",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100001",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100011",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100100",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001100110",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101000",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101001",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101011",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101101",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001101110",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110000",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110010",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110011",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110101",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001110110",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111000",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111010",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111011",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111101",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110001111111",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000000",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000010",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000100",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000101",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010000111",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001000",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001010",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001100",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001101",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010001111",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010001",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010010",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010100",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010110",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010010111",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011001",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011011",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011100",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011110",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010011111",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100001",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100011",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100100",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010100110",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101000",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101001",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101011",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101101",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010101110",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110000",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110001",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110011",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110101",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010110110",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111000",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111010",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111011",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111101",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110010111111",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000000",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000010",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000011",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000101",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011000111",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001000",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001010",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001100",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001101",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011001111",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010001",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010010",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010100",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010101",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011010111",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011001",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011010",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011100",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011110",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011011111",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100001",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100011",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100100",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011100110",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101000",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101001",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101011",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101100",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011101110",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110000",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110001",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110011",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110101",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011110110",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111000",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111010",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111011",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111101",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110011111110",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000000",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000010",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000011",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000101",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100000111",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001000",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001010",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001100",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001101",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100001111",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010000",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010010",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010100",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010101",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100010111",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011001",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011010",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011100",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011110",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100011111",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100001",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100010",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100100",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100110",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100100111",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101001",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101011",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101100",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100101110",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110000",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110001",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110011",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110101",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100110110",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111000",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111001",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111011",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111101",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110100111110",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000000",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000010",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000011",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000101",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101000111",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001000",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001010",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001011",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001101",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101001111",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010000",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010010",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010100",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010101",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101010111",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011001",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011010",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011100",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011101",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101011111",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100001",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100010",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100100",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100110",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101100111",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101001",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101011",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101100",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101101110",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110000",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110001",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110011",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110100",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101110110",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111000",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111001",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111011",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111101",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110101111110",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000000",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000010",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000011",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000101",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110000110",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001000",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001010",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001011",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001101",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110001111",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010000",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010010",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010100",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010101",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110010111",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011000",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011010",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011100",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011101",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110011111",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100001",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100010",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100100",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100110",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110100111",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101001",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101010",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101100",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101110",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110101111",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110001",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110011",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110100",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110110110",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111000",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111001",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111011",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111101",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110110111110",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000000",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000001",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000011",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000101",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111000110",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001000",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001010",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001011",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001101",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111001111",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010000",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010010",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010011",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010101",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111010111",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011000",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011010",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011100",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011101",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111011111",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100001",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100010",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100100",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100101",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111100111",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101001",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101010",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101100",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101110",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111101111",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110001",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110011",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110100",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110110",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111110111",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111001",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111011",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111100",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100110111111110",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000000",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000001",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000011",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000101",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000000110",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001000",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001010",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001011",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001101",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000001110",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010000",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010010",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010011",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010101",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000010111",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011000",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011010",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011100",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011101",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000011111",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100000",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100010",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100100",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100101",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000100111",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101001",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101010",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101100",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101110",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000101111",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110001",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110010",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110100",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110110",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000110111",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111001",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111011",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111100",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111000111110",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000000",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000001",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000011",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000100",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001000110",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001000",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001001",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001011",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001101",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001001110",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010000",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010010",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010011",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010101",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001010111",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011000",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011010",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011011",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011101",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001011111",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100000",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100010",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100100",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100101",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001100111",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101001",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101010",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101100",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101101",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001101111",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110001",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110010",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110100",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110110",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001110111",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111001",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111011",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111100",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111110",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111001111111",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000001",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000011",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000100",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010000110",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001000",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001001",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001011",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001101",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010001110",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010000",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010001",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010011",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010101",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010010110",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011000",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011010",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011011",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011101",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010011111",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100000",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100010",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100100",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100101",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010100111",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101000",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101010",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101100",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101101",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010101111",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110001",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110010",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110100",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110110",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010110111",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111001",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111010",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111100",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111110",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111010111111",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000001",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000011",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000100",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011000110",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001000",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001001",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001011",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001100",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011001110",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010000",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010001",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010011",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010101",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011010110",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011000",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011010",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011011",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011101",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011011111",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100000",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100010",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100011",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100101",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011100111",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101000",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101010",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101100",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101101",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011101111",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110001",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110010",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110100",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110101",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011110111",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111001",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111010",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111100",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111110",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111011111111",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000001",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000011",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000100",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000110",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100000111",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001001",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001011",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001100",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100001110",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010000",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010001",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010011",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010101",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100010110",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011000",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011001",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011011",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011101",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100011110",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100000",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100010",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100011",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100101",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100100111",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101000",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101010",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101100",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101101",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100101111",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110000",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110010",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110100",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110101",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100110111",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111001",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111010",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111100",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111110",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111100111111",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000001",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000010",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000100",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000110",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101000111",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001001",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001011",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001100",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101001110",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010000",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010001",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010011",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010100",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101010110",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011000",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011001",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011011",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011101",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101011110",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100000",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100010",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100011",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100101",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101100110",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101000",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101010",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101011",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101101",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101101111",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110000",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110010",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110100",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110101",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101110111",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111001",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111010",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111100",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111101",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111101111111",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000001",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000010",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000100",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000110",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110000111",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001001",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001011",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001100",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001110",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110001111",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010001",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010011",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010100",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110010110",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011000",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011001",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011011",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011101",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110011110",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100000",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100001",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100011",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100101",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110100110",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101000",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101010",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101011",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101101",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110101111",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110000",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110010",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110011",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110101",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110110111",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111000",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111010",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111100",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111101",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111110111111",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000001",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000010",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000100",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000110",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111000111",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001001",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001010",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001100",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001110",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111001111",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010001",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010011",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010100",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111010110",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011000",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011001",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011011",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011100",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111011110",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100000",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100001",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100011",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100101",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111100110",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101000",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101010",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101011",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101101",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111101110",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110000",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110010",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110011",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110101",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111110111",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111000",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111010",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111100",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111101",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1100111111111111",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000001",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000010",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000100",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000101",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000000111",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001001",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001010",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001100",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001110",
"1101000000001111",
"1101000000001111",
"1101000000001111",
"1101000000001111",
"1101000000001111",
"1101000000001111",
"1101000000001111"
);
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "block";
begin
    --ROM process
    process(clk)
    begin
        if clk'event and clk = '1' then
            data <= ROM(conv_integer(addr));
        end if;
    end process;

end Behavioral;
