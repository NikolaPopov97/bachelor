----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 09/17/2022 04:16:05 PM
-- Design Name: 
-- Module Name: phaser_datapath_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.all;
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

use STD.textio.all;
use ieee.std_logic_textio.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity phaser_datapath_tb is
--  Port ( );
end phaser_datapath_tb;

architecture Behavioral of phaser_datapath_tb is
    constant half_period: time := 10ns;
    signal on_in_s : STD_LOGIC;
    signal clk :  STD_LOGIC := '0';
    signal input_in_s : STD_LOGIC_VECTOR (15 downto 0) := x"0000";
    signal output_out_s : SIGNED(15 downto 0);
    signal reset : std_logic;
    signal out_valid: std_logic;
    type audio_type is array (104590 downto 0) of std_logic_vector(15 downto 0);
    
    signal AUDIO : audio_type :=
    ("1111111111111000",
    "1111111111111100",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111110111",
    "1111111111111001",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111101110",
    "1111111111101110",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110101",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101110",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111101111",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111101111",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111101111",
    "1111111111110000",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101111",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111110111",
    "1111111111110101",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111111",
    "1111111111111111",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101100",
    "1111111111101011",
    "1111111111101011",
    "1111111111101100",
    "1111111111101110",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111110111",
    "1111111111110011",
    "1111111111101110",
    "1111111111101010",
    "1111111111100111",
    "1111111111100110",
    "1111111111101000",
    "1111111111101010",
    "1111111111101101",
    "1111111111110000",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111001",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111101101",
    "1111111111101011",
    "1111111111101011",
    "1111111111101101",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110101",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111110000",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110100",
    "1111111111110010",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111100",
    "1111111111111010",
    "1111111111110110",
    "1111111111110011",
    "1111111111110000",
    "1111111111101111",
    "1111111111101111",
    "1111111111110000",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111110110",
    "1111111111110011",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110111",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110101",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110101",
    "1111111111110001",
    "1111111111101101",
    "1111111111101010",
    "1111111111100111",
    "1111111111100110",
    "1111111111100111",
    "1111111111101001",
    "1111111111101100",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110101",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111110110",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111000",
    "1111111111110101",
    "1111111111110010",
    "1111111111110000",
    "1111111111101111",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110111",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111010",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110111",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110010",
    "1111111111110010",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110101",
    "1111111111110101",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110101",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111101110",
    "1111111111110000",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111011",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111011",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111011",
    "1111111111111100",
    "1111111111110110",
    "1111111111110000",
    "1111111111101100",
    "1111111111101011",
    "1111111111101100",
    "1111111111101111",
    "1111111111110100",
    "1111111111111010",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110101",
    "1111111111110111",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111010",
    "1111111111111110",
    "1111111111111011",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110100",
    "1111111111111001",
    "1111111111111111",
    "1111111111111001",
    "1111111111110011",
    "1111111111101111",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110101",
    "1111111111110011",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110000",
    "1111111111101101",
    "1111111111101011",
    "1111111111101010",
    "1111111111101010",
    "1111111111101011",
    "1111111111101110",
    "1111111111110001",
    "1111111111110101",
    "1111111111111001",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110011",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101110",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000",
    "1111111111110011",
    "1111111111110000",
    "1111111111101110",
    "1111111111101110",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111111011",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111011",
    "1111111111111101",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111010",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110101",
    "1111111111110011",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111111001",
    "1111111111111101",
    "1111111111111011",
    "1111111111110110",
    "1111111111110010",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110111",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110111",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110111",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111110111",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111100",
    "1111111111111101",
    "1111111111111000",
    "1111111111110011",
    "1111111111110000",
    "1111111111101111",
    "1111111111110000",
    "1111111111110011",
    "1111111111110111",
    "1111111111111011",
    "1111111111111111",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110111",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111011",
    "1111111111111111",
    "1111111111111010",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110101",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111010",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110101",
    "1111111111110111",
    "1111111111111011",
    "1111111111111101",
    "1111111111111000",
    "1111111111110011",
    "1111111111101110",
    "1111111111101100",
    "1111111111101100",
    "1111111111101111",
    "1111111111110011",
    "1111111111111001",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000",
    "1111111111110101",
    "1111111111110011",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111010",
    "1111111111111101",
    "1111111111111011",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101011",
    "1111111111101100",
    "1111111111101110",
    "1111111111110011",
    "1111111111110110",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110101",
    "1111111111110011",
    "1111111111110000",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110010",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111101111",
    "1111111111101010",
    "1111111111100110",
    "1111111111100011",
    "1111111111100010",
    "1111111111100011",
    "1111111111100101",
    "1111111111101000",
    "1111111111101101",
    "1111111111110011",
    "1111111111111001",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110110",
    "1111111111111011",
    "1111111111111100",
    "1111111111110110",
    "1111111111110001",
    "1111111111101110",
    "1111111111101101",
    "1111111111101110",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111111",
    "1111111111111010",
    "1111111111110101",
    "1111111111110000",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101110",
    "1111111111110001",
    "1111111111110101",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111101110",
    "1111111111101111",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111101111",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110011",
    "1111111111110110",
    "1111111111111011",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110010",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110100",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111111000",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110111",
    "1111111111111010",
    "1111111111111100",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111101111",
    "1111111111101110",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111010",
    "1111111111110110",
    "1111111111110011",
    "1111111111110010",
    "1111111111110011",
    "1111111111110101",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111111",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111011",
    "1111111111111101",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111001",
    "1111111111110100",
    "1111111111101111",
    "1111111111101011",
    "1111111111101001",
    "1111111111101001",
    "1111111111101100",
    "1111111111110000",
    "1111111111110101",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111111",
    "1111111111111101",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110000",
    "1111111111101101",
    "1111111111101011",
    "1111111111101100",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111110110",
    "1111111111110011",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110101",
    "1111111111110010",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110000",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111010",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110101",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110011",
    "1111111111101110",
    "1111111111101000",
    "1111111111100011",
    "1111111111011110",
    "1111111111011011",
    "1111111111011010",
    "1111111111011100",
    "1111111111100001",
    "1111111111101000",
    "1111111111110011",
    "1111111111111110",
    "1111111111110011",
    "1111111111100111",
    "1111111111011110",
    "1111111111010110",
    "1111111111010001",
    "1111111111001111",
    "1111111111010001",
    "1111111111010110",
    "1111111111011101",
    "1111111111100101",
    "1111111111101110",
    "1111111111110111",
    "1111111111111110",
    "1111111111111000",
    "1111111111110011",
    "1111111111110000",
    "1111111111101111",
    "1111111111110000",
    "1111111111110011",
    "1111111111111000",
    "1111111111111101",
    "1111111111111010",
    "1111111111110101",
    "1111111111110001",
    "1111111111101110",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111111",
    "1111111111111111",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111101111",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110100",
    "1111111111110110",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111110110",
    "1111111111101111",
    "1111111111100111",
    "1111111111100000",
    "1111111111011000",
    "1111111111010010",
    "1111111111001101",
    "1111111111001011",
    "1111111111001100",
    "1111111111010000",
    "1111111111011000",
    "1111111111100011",
    "1111111111110000",
    "1111111111111101",
    "1111111111101110",
    "1111111111100010",
    "1111111111010111",
    "1111111111010001",
    "1111111111001111",
    "1111111111010010",
    "1111111111011010",
    "1111111111100101",
    "1111111111110010",
    "1111111111111101",
    "1111111111110000",
    "1111111111100110",
    "1111111111011111",
    "1111111111011011",
    "1111111111011010",
    "1111111111011100",
    "1111111111011111",
    "1111111111100011",
    "1111111111101001",
    "1111111111101110",
    "1111111111110011",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110101",
    "1111111111110011",
    "1111111111110000",
    "1111111111101101",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110101",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111010",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000",
    "1111111111110010",
    "1111111111101011",
    "1111111111100110",
    "1111111111100001",
    "1111111111011110",
    "1111111111011100",
    "1111111111011100",
    "1111111111011111",
    "1111111111100100",
    "1111111111101101",
    "1111111111111001",
    "1111111111111000",
    "1111111111101010",
    "1111111111011111",
    "1111111111010111",
    "1111111111010001",
    "1111111111001111",
    "1111111111010000",
    "1111111111010101",
    "1111111111011100",
    "1111111111100100",
    "1111111111101110",
    "1111111111111000",
    "1111111111111101",
    "1111111111110110",
    "1111111111110010",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111010",
    "1111111111111111",
    "1111111111111001",
    "1111111111110100",
    "1111111111110000",
    "1111111111101100",
    "1111111111101010",
    "1111111111101010",
    "1111111111101011",
    "1111111111101110",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110000",
    "1111111111101100",
    "1111111111101010",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111110000",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111000",
    "1111111111110101",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111111001",
    "1111111111111011",
    "1111111111111111",
    "1111111111111011",
    "1111111111110110",
    "1111111111110001",
    "1111111111101110",
    "1111111111101100",
    "1111111111101100",
    "1111111111101101",
    "1111111111110000",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111110",
    "1111111111111001",
    "1111111111110011",
    "1111111111101011",
    "1111111111100100",
    "1111111111011110",
    "1111111111011001",
    "1111111111010110",
    "1111111111010101",
    "1111111111011000",
    "1111111111011111",
    "1111111111101000",
    "1111111111110101",
    "1111111111111011",
    "1111111111101110",
    "1111111111100100",
    "1111111111011110",
    "1111111111011011",
    "1111111111011011",
    "1111111111011110",
    "1111111111100010",
    "1111111111101000",
    "1111111111110000",
    "1111111111110111",
    "1111111111111111",
    "1111111111111000",
    "1111111111110011",
    "1111111111101110",
    "1111111111101011",
    "1111111111101010",
    "1111111111101001",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111101110",
    "1111111111110010",
    "1111111111110111",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110001",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101100",
    "1111111111101011",
    "1111111111101100",
    "1111111111110000",
    "1111111111110011",
    "1111111111111000",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111110",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111110110",
    "1111111111110011",
    "1111111111101111",
    "1111111111101011",
    "1111111111101000",
    "1111111111100101",
    "1111111111100010",
    "1111111111100000",
    "1111111111011101",
    "1111111111011100",
    "1111111111011101",
    "1111111111100001",
    "1111111111100110",
    "1111111111101100",
    "1111111111110011",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111110110",
    "1111111111110000",
    "1111111111100110",
    "1111111111011101",
    "1111111111010100",
    "1111111111001100",
    "1111111111000110",
    "1111111111000011",
    "1111111111000010",
    "1111111111000100",
    "1111111111001001",
    "1111111111010000",
    "1111111111011011",
    "1111111111100110",
    "1111111111110011",
    "1111111111111111",
    "1111111111110100",
    "1111111111101011",
    "1111111111100101",
    "1111111111100010",
    "1111111111100011",
    "1111111111100110",
    "1111111111101100",
    "1111111111110011",
    "1111111111111100",
    "1111111111111001",
    "1111111111110001",
    "1111111111101011",
    "1111111111100110",
    "1111111111100100",
    "1111111111100011",
    "1111111111100101",
    "1111111111100111",
    "1111111111101010",
    "1111111111101110",
    "1111111111110011",
    "1111111111111000",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101110",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111010",
    "1111111111110111",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110111",
    "1111111111111010",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111101110",
    "1111111111101110",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110100",
    "1111111111111000",
    "1111111111111100",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111010",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110010",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110101",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111110101",
    "1111111111110000",
    "1111111111101010",
    "1111111111100101",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100100",
    "1111111111100111",
    "1111111111101011",
    "1111111111110000",
    "1111111111110110",
    "1111111111111111",
    "1111111111110100",
    "1111111111101001",
    "1111111111011111",
    "1111111111010111",
    "1111111111010010",
    "1111111111010001",
    "1111111111010011",
    "1111111111011000",
    "1111111111011100",
    "1111111111100000",
    "1111111111100010",
    "1111111111100100",
    "1111111111100110",
    "1111111111100110",
    "1111111111100100",
    "1111111111100010",
    "1111111111011100",
    "1111111111010110",
    "1111111111010000",
    "1111111111001100",
    "1111111111001100",
    "1111111111010001",
    "1111111111011100",
    "1111111111101010",
    "1111111111111101",
    "1111111111101011",
    "1111111111010110",
    "1111111111000001",
    "1111111110101111",
    "1111111110100010",
    "1111111110011001",
    "1111111110010110",
    "1111111110010111",
    "1111111110011101",
    "1111111110100101",
    "1111111110110000",
    "1111111110111101",
    "1111111111001010",
    "1111111111011001",
    "1111111111100110",
    "1111111111110000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110011",
    "1111111111101110",
    "1111111111101001",
    "1111111111100100",
    "1111111111011111",
    "1111111111011011",
    "1111111111011000",
    "1111111111010111",
    "1111111111011001",
    "1111111111011101",
    "1111111111100010",
    "1111111111100110",
    "1111111111101011",
    "1111111111101110",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111101110",
    "1111111111101100",
    "1111111111101010",
    "1111111111101000",
    "1111111111100110",
    "1111111111100101",
    "1111111111100101",
    "1111111111100101",
    "1111111111100110",
    "1111111111101000",
    "1111111111101011",
    "1111111111101101",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111101111",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101100",
    "1111111111101011",
    "1111111111101011",
    "1111111111101011",
    "1111111111101011",
    "1111111111101100",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110011",
    "1111111111110110",
    "1111111111111000",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110100",
    "1111111111101111",
    "1111111111101010",
    "1111111111100111",
    "1111111111100100",
    "1111111111100010",
    "1111111111100010",
    "1111111111100100",
    "1111111111100111",
    "1111111111101011",
    "1111111111101101",
    "1111111111101101",
    "1111111111101011",
    "1111111111101000",
    "1111111111100110",
    "1111111111100100",
    "1111111111100101",
    "1111111111101000",
    "1111111111101011",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111101111",
    "1111111111101111",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110001",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110000",
    "1111111111101101",
    "1111111111101010",
    "1111111111100110",
    "1111111111100001",
    "1111111111011011",
    "1111111111010101",
    "1111111111010000",
    "1111111111001101",
    "1111111111001101",
    "1111111111001111",
    "1111111111010100",
    "1111111111011011",
    "1111111111100011",
    "1111111111101101",
    "1111111111110110",
    "1111111111111110",
    "1111111111111001",
    "1111111111110101",
    "1111111111110011",
    "1111111111110100",
    "1111111111110111",
    "1111111111111011",
    "1111111111111111",
    "1111111111111001",
    "1111111111110101",
    "1111111111110000",
    "1111111111101011",
    "1111111111100111",
    "1111111111100011",
    "1111111111100000",
    "1111111111011101",
    "1111111111011011",
    "1111111111011001",
    "1111111111011001",
    "1111111111011011",
    "1111111111011110",
    "1111111111100010",
    "1111111111100111",
    "1111111111101101",
    "1111111111110010",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111101110",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110010",
    "1111111111110100",
    "1111111111110110",
    "1111111111111010",
    "1111111111111101",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111101110",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110100",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101110",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111001",
    "1111111111110100",
    "1111111111110000",
    "1111111111101110",
    "1111111111101100",
    "1111111111101011",
    "1111111111101011",
    "1111111111101100",
    "1111111111101101",
    "1111111111101111",
    "1111111111110001",
    "1111111111110100",
    "1111111111110111",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111111000",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111011",
    "1111111111111111",
    "1111111111111010",
    "1111111111110101",
    "1111111111110000",
    "1111111111101100",
    "1111111111101001",
    "1111111111101000",
    "1111111111100111",
    "1111111111100111",
    "1111111111101001",
    "1111111111101011",
    "1111111111101110",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111001",
    "1111111111110110",
    "1111111111110010",
    "1111111111101101",
    "1111111111101000",
    "1111111111100101",
    "1111111111100100",
    "1111111111100110",
    "1111111111101010",
    "1111111111110011",
    "1111111111111100",
    "1111111111110110",
    "1111111111101011",
    "1111111111100001",
    "1111111111011000",
    "1111111111010001",
    "1111111111001111",
    "1111111111010001",
    "1111111111011000",
    "1111111111100001",
    "1111111111101101",
    "1111111111111010",
    "1111111111110110",
    "1111111111101010",
    "1111111111100010",
    "1111111111011011",
    "1111111111010110",
    "1111111111010101",
    "1111111111010101",
    "1111111111011000",
    "1111111111011101",
    "1111111111100100",
    "1111111111101101",
    "1111111111110110",
    "1111111111111110",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101101",
    "1111111111110000",
    "1111111111110011",
    "1111111111111001",
    "1111111111111100",
    "1111111111110101",
    "1111111111101110",
    "1111111111101000",
    "1111111111100100",
    "1111111111100011",
    "1111111111100100",
    "1111111111101000",
    "1111111111101111",
    "1111111111111000",
    "1111111111111101",
    "1111111111110110",
    "1111111111110000",
    "1111111111101110",
    "1111111111110000",
    "1111111111110110",
    "1111111111111110",
    "1111111111110011",
    "1111111111100110",
    "1111111111011100",
    "1111111111010101",
    "1111111111010001",
    "1111111111010010",
    "1111111111010110",
    "1111111111011101",
    "1111111111100110",
    "1111111111101111",
    "1111111111111000",
    "1111111111111100",
    "1111111111110011",
    "1111111111101011",
    "1111111111100011",
    "1111111111011100",
    "1111111111010111",
    "1111111111010011",
    "1111111111010000",
    "1111111111001111",
    "1111111111001110",
    "1111111111001100",
    "1111111111001010",
    "1111111111001000",
    "1111111111000110",
    "1111111111000100",
    "1111111111000011",
    "1111111111000011",
    "1111111111000101",
    "1111111111000110",
    "1111111111001001",
    "1111111111001101",
    "1111111111010010",
    "1111111111011000",
    "1111111111011111",
    "1111111111101000",
    "1111111111110010",
    "1111111111111101",
    "1111111111110011",
    "1111111111101000",
    "1111111111011110",
    "1111111111010101",
    "1111111111001111",
    "1111111111001011",
    "1111111111001010",
    "1111111111001011",
    "1111111111001101",
    "1111111111010000",
    "1111111111010011",
    "1111111111010111",
    "1111111111011011",
    "1111111111011110",
    "1111111111100001",
    "1111111111100011",
    "1111111111100101",
    "1111111111100110",
    "1111111111101000",
    "1111111111101010",
    "1111111111101100",
    "1111111111101111",
    "1111111111110001",
    "1111111111110010",
    "1111111111110001",
    "1111111111110000",
    "1111111111101110",
    "1111111111101100",
    "1111111111101010",
    "1111111111101000",
    "1111111111100111",
    "1111111111100110",
    "1111111111100101",
    "1111111111100100",
    "1111111111100100",
    "1111111111100101",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101011",
    "1111111111101010",
    "1111111111101001",
    "1111111111100110",
    "1111111111100100",
    "1111111111100011",
    "1111111111100011",
    "1111111111100101",
    "1111111111100111",
    "1111111111101010",
    "1111111111101100",
    "1111111111101100",
    "1111111111101010",
    "1111111111100110",
    "1111111111100010",
    "1111111111011101",
    "1111111111011000",
    "1111111111010101",
    "1111111111010100",
    "1111111111010110",
    "1111111111011010",
    "1111111111100000",
    "1111111111100111",
    "1111111111110000",
    "1111111111111010",
    "1111111111111001",
    "1111111111110000",
    "1111111111101000",
    "1111111111100011",
    "1111111111100000",
    "1111111111011111",
    "1111111111100000",
    "1111111111100100",
    "1111111111101100",
    "1111111111110110",
    "1111111111111001",
    "1111111111101011",
    "1111111111011100",
    "1111111111001101",
    "1111111111000010",
    "1111111110111010",
    "1111111110110101",
    "1111111110110110",
    "1111111110111011",
    "1111111111000011",
    "1111111111001101",
    "1111111111011011",
    "1111111111101001",
    "1111111111111000",
    "1111111111111000",
    "1111111111101101",
    "1111111111100101",
    "1111111111100010",
    "1111111111100011",
    "1111111111100111",
    "1111111111101100",
    "1111111111110001",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111011",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110000",
    "1111111111101111",
    "1111111111101111",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110110",
    "1111111111110110",
    "1111111111110111",
    "1111111111110111",
    "1111111111110111",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111101111",
    "1111111111101110",
    "1111111111101100",
    "1111111111101001",
    "1111111111100101",
    "1111111111100010",
    "1111111111011111",
    "1111111111011101",
    "1111111111011100",
    "1111111111011100",
    "1111111111011100",
    "1111111111011100",
    "1111111111011011",
    "1111111111011001",
    "1111111111011001",
    "1111111111011001",
    "1111111111011010",
    "1111111111011100",
    "1111111111011111",
    "1111111111100001",
    "1111111111100011",
    "1111111111100100",
    "1111111111100101",
    "1111111111100111",
    "1111111111101010",
    "1111111111101100",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110001",
    "1111111111101110",
    "1111111111101100",
    "1111111111101011",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101001",
    "1111111111101000",
    "1111111111100111",
    "1111111111100110",
    "1111111111100100",
    "1111111111100011",
    "1111111111100011",
    "1111111111100011",
    "1111111111100101",
    "1111111111101000",
    "1111111111101100",
    "1111111111110000",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111101111",
    "1111111111101001",
    "1111111111100010",
    "1111111111011010",
    "1111111111010001",
    "1111111111001010",
    "1111111111000110",
    "1111111111000100",
    "1111111111000111",
    "1111111111001101",
    "1111111111010111",
    "1111111111100010",
    "1111111111101101",
    "1111111111111001",
    "1111111111111010",
    "1111111111110011",
    "1111111111101101",
    "1111111111101010",
    "1111111111101011",
    "1111111111101110",
    "1111111111110011",
    "1111111111111001",
    "1111111111111100",
    "1111111111110011",
    "1111111111101100",
    "1111111111100110",
    "1111111111100010",
    "1111111111100000",
    "1111111111011111",
    "1111111111011111",
    "1111111111100000",
    "1111111111100010",
    "1111111111100011",
    "1111111111100100",
    "1111111111100101",
    "1111111111101000",
    "1111111111101011",
    "1111111111110000",
    "1111111111110100",
    "1111111111111010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111010",
    "1111111111111001",
    "1111111111111001",
    "1111111111110111",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110010",
    "1111111111110001",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111101101",
    "1111111111101011",
    "1111111111101001",
    "1111111111101000",
    "1111111111101000",
    "1111111111101000",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111101101",
    "1111111111101110",
    "1111111111101110",
    "1111111111101110",
    "1111111111101101",
    "1111111111101100",
    "1111111111101100",
    "1111111111101011",
    "1111111111101011",
    "1111111111101011",
    "1111111111101010",
    "1111111111101010",
    "1111111111101001",
    "1111111111101001",
    "1111111111101001",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101010",
    "1111111111101000",
    "1111111111100111",
    "1111111111100110",
    "1111111111100110",
    "1111111111101000",
    "1111111111101100",
    "1111111111110001",
    "1111111111110111",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111110111",
    "1111111111110011",
    "1111111111101110",
    "1111111111101100",
    "1111111111101100",
    "1111111111101110",
    "1111111111110011",
    "1111111111111001",
    "1111111111111100",
    "1111111111110100",
    "1111111111101101",
    "1111111111100111",
    "1111111111100011",
    "1111111111100011",
    "1111111111100111",
    "1111111111101101",
    "1111111111110111",
    "1111111111111011",
    "1111111111101111",
    "1111111111100100",
    "1111111111011100",
    "1111111111010110",
    "1111111111010001",
    "1111111111010000",
    "1111111111001111",
    "1111111111001111",
    "1111111111010000",
    "1111111111010001",
    "1111111111010010",
    "1111111111010110",
    "1111111111011011",
    "1111111111100010",
    "1111111111101001",
    "1111111111110000",
    "1111111111111000",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111100",
    "1111111111111011",
    "1111111111111000",
    "1111111111110011",
    "1111111111101100",
    "1111111111100011",
    "1111111111010111",
    "1111111111001001",
    "1111111110111100",
    "1111111110101111",
    "1111111110100101",
    "1111111110100001",
    "1111111110100010",
    "1111111110101001",
    "1111111110110111",
    "1111111111001000",
    "1111111111011101",
    "1111111111110011",
    "1111111111110110",
    "1111111111100010",
    "1111111111010000",
    "1111111111000001",
    "1111111110110101",
    "1111111110101100",
    "1111111110101000",
    "1111111110100110",
    "1111111110101000",
    "1111111110101100",
    "1111111110110010",
    "1111111110111010",
    "1111111111000011",
    "1111111111001011",
    "1111111111010100",
    "1111111111011100",
    "1111111111100010",
    "1111111111100110",
    "1111111111100111",
    "1111111111100111",
    "1111111111100101",
    "1111111111100010",
    "1111111111011110",
    "1111111111011011",
    "1111111111011001",
    "1111111111011001",
    "1111111111011001",
    "1111111111011011",
    "1111111111011110",
    "1111111111100001",
    "1111111111100100",
    "1111111111100111",
    "1111111111101001",
    "1111111111101010",
    "1111111111101010",
    "1111111111101001",
    "1111111111100111",
    "1111111111100100",
    "1111111111100001",
    "1111111111011101",
    "1111111111011001",
    "1111111111010110",
    "1111111111010100",
    "1111111111010010",
    "1111111111010010",
    "1111111111010100",
    "1111111111010110",
    "1111111111011000",
    "1111111111011001",
    "1111111111011010",
    "1111111111011011",
    "1111111111011011",
    "1111111111011011",
    "1111111111011011",
    "1111111111011100",
    "1111111111011101",
    "1111111111011111",
    "1111111111100001",
    "1111111111100010",
    "1111111111100100",
    "1111111111100110",
    "1111111111101000",
    "1111111111101000",
    "1111111111101000",
    "1111111111101000",
    "1111111111100111",
    "1111111111100111",
    "1111111111101000",
    "1111111111101001",
    "1111111111101100",
    "1111111111101110",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111101111",
    "1111111111101101",
    "1111111111101011",
    "1111111111101010",
    "1111111111101011",
    "1111111111101101",
    "1111111111110001",
    "1111111111110110",
    "1111111111111011",
    "1111111111111101",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111101101",
    "1111111111101011",
    "1111111111101001",
    "1111111111100111",
    "1111111111100110",
    "1111111111100100",
    "1111111111100011",
    "1111111111100011",
    "1111111111100011",
    "1111111111100100",
    "1111111111100110",
    "1111111111101010",
    "1111111111101101",
    "1111111111110001",
    "1111111111110011",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110001",
    "1111111111110000",
    "1111111111101111",
    "1111111111101110",
    "1111111111101101",
    "1111111111101100",
    "1111111111101010",
    "1111111111100111",
    "1111111111100011",
    "1111111111011110",
    "1111111111011001",
    "1111111111010101",
    "1111111111010001",
    "1111111111010000",
    "1111111111010001",
    "1111111111010101",
    "1111111111011010",
    "1111111111100000",
    "1111111111100100",
    "1111111111100111",
    "1111111111100111",
    "1111111111100101",
    "1111111111011111",
    "1111111111010111",
    "1111111111001101",
    "1111111111000011",
    "1111111110111001",
    "1111111110101111",
    "1111111110101001",
    "1111111110100111",
    "1111111110101001",
    "1111111110101110",
    "1111111110110110",
    "1111111111000010",
    "1111111111001101",
    "1111111111011001",
    "1111111111100100",
    "1111111111101101",
    "1111111111110101",
    "1111111111111010",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111101110",
    "1111111111100111",
    "1111111111100001",
    "1111111111011010",
    "1111111111010011",
    "1111111111001110",
    "1111111111001010",
    "1111111111001001",
    "1111111111001001",
    "1111111111001100",
    "1111111111001111",
    "1111111111010100",
    "1111111111011001",
    "1111111111011101",
    "1111111111100001",
    "1111111111100010",
    "1111111111100011",
    "1111111111100011",
    "1111111111100001",
    "1111111111011110",
    "1111111111011100",
    "1111111111011001",
    "1111111111011001",
    "1111111111011010",
    "1111111111011101",
    "1111111111100001",
    "1111111111100101",
    "1111111111101000",
    "1111111111101001",
    "1111111111101001",
    "1111111111101000",
    "1111111111101000",
    "1111111111101000",
    "1111111111101010",
    "1111111111101100",
    "1111111111101110",
    "1111111111110001",
    "1111111111110011",
    "1111111111110100",
    "1111111111110100",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110000",
    "1111111111101110",
    "1111111111101100",
    "1111111111101011",
    "1111111111101011",
    "1111111111101011",
    "1111111111101101",
    "1111111111110000",
    "1111111111110011",
    "1111111111110110",
    "1111111111111010",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110010",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110100",
    "1111111111110011",
    "1111111111110010",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110001",
    "1111111111110010",
    "1111111111110011",
    "1111111111110011",
    "1111111111110100",
    "1111111111110101",
    "1111111111110110",
    "1111111111110110",
    "1111111111111000",
    "1111111111111001",
    "1111111111111001",
    "1111111111111011",
    "1111111111111011",
    "1111111111111001",
    "1111111111110110",
    "1111111111110001",
    "1111111111101011",
    "1111111111100100",
    "1111111111011111",
    "1111111111011011",
    "1111111111011010",
    "1111111111011010",
    "1111111111011101",
    "1111111111100010",
    "1111111111100111",
    "1111111111101101",
    "1111111111110100",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111110110",
    "1111111111110000",
    "1111111111101001",
    "1111111111100011",
    "1111111111011110",
    "1111111111011010",
    "1111111111011000",
    "1111111111011000",
    "1111111111011100",
    "1111111111100010",
    "1111111111101010",
    "1111111111110100",
    "1111111111111110",
    "1111111111110110",
    "1111111111101110",
    "1111111111101010",
    "1111111111101001",
    "1111111111101011",
    "1111111111110000",
    "1111111111110110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110000",
    "1111111111101000",
    "1111111111100000",
    "1111111111011001",
    "1111111111010011",
    "1111111111001111",
    "1111111111001101",
    "1111111111001101",
    "1111111111001111",
    "1111111111010010",
    "1111111111010101",
    "1111111111011000",
    "1111111111011011",
    "1111111111011110",
    "1111111111100001",
    "1111111111100100",
    "1111111111100111",
    "1111111111101011",
    "1111111111110000",
    "1111111111110100",
    "1111111111111011",
    "1111111111111100",
    "1111111111110111",
    "1111111111110011",
    "1111111111110000",
    "1111111111110000",
    "1111111111110001",
    "1111111111110100",
    "1111111111111001",
    "1111111111111101",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110001",
    "1111111111101110",
    "1111111111101100",
    "1111111111101010",
    "1111111111101000",
    "1111111111100110",
    "1111111111100100",
    "1111111111100010",
    "1111111111100001",
    "1111111111011110",
    "1111111111011011",
    "1111111111011000",
    "1111111111010110",
    "1111111111010100",
    "1111111111010011",
    "1111111111010010",
    "1111111111010010",
    "1111111111010010",
    "1111111111010011",
    "1111111111010110",
    "1111111111011001",
    "1111111111011110",
    "1111111111100100",
    "1111111111101011",
    "1111111111110100",
    "1111111111111101",
    "1111111111110110",
    "1111111111101100",
    "1111111111100011",
    "1111111111011011",
    "1111111111010010",
    "1111111111001011",
    "1111111111000111",
    "1111111111000100",
    "1111111111000100",
    "1111111111000110",
    "1111111111001010",
    "1111111111001111",
    "1111111111010110",
    "1111111111011101",
    "1111111111100100",
    "1111111111101011",
    "1111111111110011",
    "1111111111111010",
    "1111111111111011",
    "1111111111110010",
    "1111111111101001",
    "1111111111100011",
    "1111111111011110",
    "1111111111011100",
    "1111111111011011",
    "1111111111011100",
    "1111111111011101",
    "1111111111011110",
    "1111111111011111",
    "1111111111011111",
    "1111111111011110",
    "1111111111011101",
    "1111111111011101",
    "1111111111011100",
    "1111111111011100",
    "1111111111011110",
    "1111111111100000",
    "1111111111100100",
    "1111111111101001",
    "1111111111110000",
    "1111111111110110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111110110",
    "1111111111110100",
    "1111111111110011",
    "1111111111110000",
    "1111111111101110",
    "1111111111101011",
    "1111111111101010",
    "1111111111101001",
    "1111111111101001",
    "1111111111101010",
    "1111111111101100",
    "1111111111110000",
    "1111111111110100",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111111000",
    "1111111111111001",
    "1111111111111101",
    "1111111111111011",
    "1111111111110100",
    "1111111111101111",
    "1111111111101011",
    "1111111111101001",
    "1111111111101011",
    "1111111111110000",
    "1111111111111001",
    "1111111111111010",
    "1111111111101110",
    "1111111111100010",
    "1111111111010111",
    "1111111111001110",
    "1111111111001001",
    "1111111111001000",
    "1111111111001011",
    "1111111111010001",
    "1111111111011001",
    "1111111111100010",
    "1111111111101100",
    "1111111111110111",
    "1111111111111100",
    "1111111111110001",
    "1111111111100110",
    "1111111111011110",
    "1111111111011000",
    "1111111111010110",
    "1111111111011000",
    "1111111111011101",
    "1111111111100011",
    "1111111111101011",
    "1111111111110011",
    "1111111111111001",
    "1111111111111111",
    "1111111111111010",
    "1111111111110110",
    "1111111111110010",
    "1111111111110000",
    "1111111111101101",
    "1111111111101101",
    "1111111111101101",
    "1111111111101110",
    "1111111111101111",
    "1111111111101110",
    "1111111111101100",
    "1111111111101010",
    "1111111111100111",
    "1111111111100101",
    "1111111111100100",
    "1111111111100100",
    "1111111111100101",
    "1111111111101000",
    "1111111111101100",
    "1111111111110000",
    "1111111111110101",
    "1111111111111001",
    "1111111111111011",
    "1111111111111100",
    "1111111111111101",
    "1111111111111111",
    "1111111111111100",
    "1111111111111001",
    "1111111111110101",
    "1111111111110000",
    "1111111111101100",
    "1111111111101001",
    "1111111111100111",
    "1111111111100110",
    "1111111111100111",
    "1111111111101001",
    "1111111111101100",
    "1111111111110001",
    "1111111111111001",
    "1111111111111101",
    "1111111111110101",
    "1111111111101110",
    "1111111111101001",
    "1111111111100111",
    "1111111111101000",
    "1111111111101100",
    "1111111111110011",
    "1111111111111010",
    "1111111111111100",
    "1111111111110110",
    "1111111111110010",
    "1111111111101111",
    "1111111111101110",
    "1111111111101110",
    "1111111111101111",
    "1111111111110001",
    "1111111111110011",
    "1111111111110111",
    "1111111111111100",
    "1111111111111100",
    "1111111111110110",
    "1111111111110001",
    "1111111111101101",
    "1111111111101001",
    "1111111111100101",
    "1111111111100010",
    "1111111111100001",
    "1111111111100001",
    "1111111111100010",
    "1111111111100110",
    "1111111111101101",
    "1111111111110101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111001",
    "1111111111111011",
    "1111111111111101",
    "1111111111110110",
    "1111111111101110",
    "1111111111100110",
    "1111111111011111",
    "1111111111011000",
    "1111111111010011",
    "1111111111010001",
    "1111111111010000",
    "1111111111010000",
    "1111111111010010",
    "1111111111010100",
    "1111111111010110",
    "1111111111010110",
    "1111111111010110",
    "1111111111010100",
    "1111111111010010",
    "1111111111010000",
    "1111111111001111",
    "1111111111001111",
    "1111111111010010",
    "1111111111010111",
    "1111111111011110",
    "1111111111100100",
    "1111111111101100",
    "1111111111110010",
    "1111111111110110",
    "1111111111111001",
    "1111111111111001",
    "1111111111111000",
    "1111111111110101",
    "1111111111110001",
    "1111111111101101",
    "1111111111101001",
    "1111111111100111",
    "1111111111100110",
    "1111111111100111",
    "1111111111101001",
    "1111111111101100",
    "1111111111110000",
    "1111111111110101",
    "1111111111111010",
    "1111111111111110",
    "1111111111111100",
    "1111111111111100",
    "1111111111111101",
    "1111111111111011",
    "1111111111110010",
    "1111111111100111",
    "1111111111011010",
    "1111111111001101",
    "1111111111000001",
    "1111111110111000",
    "1111111110110011",
    "1111111110110010",
    "1111111110110110",
    "1111111110111111",
    "1111111111001010",
    "1111111111011000",
    "1111111111100111",
    "1111111111110110",
    "1111111111111011",
    "1111111111110001",
    "1111111111101011",
    "1111111111101001",
    "1111111111101010",
    "1111111111101101",
    "1111111111110001",
    "1111111111110100",
    "1111111111111000",
    "1111111111111011",
    "1111111111111101",
    "1111111111111101",
    "1111111111111100",
    "1111111111111100",
    "1111111111111100",
    "1111111111111111",
    "1111111111111100",
    "1111111111111011",
    "1111111111111010",
    "1111111111111011",
    "1111111111111101",
    "1111111111111100",
    "1111111111110111",
    "1111111111110011",
    "1111111111101111",
    "1111111111101100",
    "1111111111101011",
    "1111111111101100",
    "1111111111101101",
    "1111111111110000",
    "1111111111110101",
    "1111111111111001",
    "1111111111111101",
    "1111111111111100",
    "1111111111111010",
    "1111111111111001",
    "1111111111111010",
    "1111111111111011",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110011",
    "1111111111101110",
    "1111111111101010",
    "1111111111100110",
    "1111111111100100",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100100",
    "1111111111100111",
    "1111111111101011",
    "1111111111110000",
    "1111111111110101",
    "1111111111111010",
    "1111111111111101",
    "1111111111111111",
    "1111111111111110",
    "1111111111111100",
    "1111111111111000",
    "1111111111110100",
    "1111111111110001",
    "1111111111101110",
    "1111111111101100",
    "1111111111101010",
    "1111111111101000",
    "1111111111100110",
    "1111111111100100",
    "1111111111100010",
    "1111111111100010",
    "1111111111100010",
    "1111111111100011",
    "1111111111100110",
    "1111111111101000",
    "1111111111101011",
    "1111111111101101",
    "1111111111101101",
    "1111111111101011",
    "1111111111100110",
    "1111111111100001",
    "1111111111011010",
    "1111111111010011",
    "1111111111001101",
    "1111111111001010",
    "1111111111001001",
    "1111111111001100",
    "1111111111010000",
    "1111111111010111",
    "1111111111011111",
    "1111111111101000",
    "1111111111110001",
    "1111111111111011",
    "1111111111111011",
    "1111111111110100",
    "1111111111110001",
    "1111111111110000",
    "1111111111110000",
    "1111111111110100",
    "1111111111111000",
    "1111111111111101",
    "1111111111111011",
    "1111111111110110",
    "1111111111110011",
    "1111111111110000",
    "1111111111101110",
    "1111111111101101",
    "1111111111101100",
    "1111111111101011",
    "1111111111101010",
    "1111111111101000",
    "1111111111100101",
    "1111111111100000",
    "1111111111011010",
    "1111111111010011",
    "1111111111001110",
    "1111111111001010",
    "1111111111001001",
    "1111111111001010",
    "1111111111001101",
    "1111111111010011",
    "1111111111011010",
    "1111111111100010",
    "1111111111101001",
    "1111111111110001",
    "1111111111111000",
    "1111111111111100",
    "1111111111111110",
    "1111111111111101",
    "1111111111111011",
    "1111111111110111",
    "1111111111110100",
    "1111111111110100",
    "1111111111111001",
    "1111111111111011",
    "1111111111101101",
    "1111111111011110",
    "1111111111001101",
    "1111111110111101",
    "1111111110101110",
    "1111111110100100",
    "1111111110011101",
    "1111111110011001",
    "1111111110011001",
    "1111111110011110",
    "1111111110100111",
    "1111111110110010",
    "1111111111000001",
    "1111111111010001",
    "1111111111100011",
    "1111111111110100",
    "1111111111111000",
    "1111111111101000",
    "1111111111011011",
    "1111111111001111",
    "1111111111000110",
    "1111111111000001",
    "1111111110111111",
    "1111111111000001",
    "1111111111000110",
    "1111111111001100",
    "1111111111010100",
    "1111111111011010",
    "1111111111011111",
    "1111111111100010",
    "1111111111100011",
    "1111111111100100",
    "1111111111100101",
    "1111111111100110",
    "1111111111100111",
    "1111111111101000",
    "1111111111101001",
    "1111111111101001",
    "1111111111101000",
    "1111111111100101",
    "1111111111100010",
    "1111111111011111",
    "1111111111011011",
    "1111111111011000",
    "1111111111010101",
    "1111111111010011",
    "1111111111010010",
    "1111111111010011",
    "1111111111010110",
    "1111111111011011",
    "1111111111100001",
    "1111111111100111",
    "1111111111101110",
    "1111111111110011",
    "1111111111110110",
    "1111111111110111",
    "1111111111110110",
    "1111111111110001",
    "1111111111101100",
    "1111111111100111",
    "1111111111100010",
    "1111111111011111",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011110",
    "1111111111011110",
    "1111111111011110",
    "1111111111011101",
    "1111111111011101",
    "1111111111011101",
    "1111111111011110",
    "1111111111011111",
    "1111111111011111",
    "1111111111100000",
    "1111111111100000",
    "1111111111100000",
    "1111111111011111",
    "1111111111011110",
    "1111111111011101",
    "1111111111011100",
    "1111111111011100",
    "1111111111011101",
    "1111111111011111",
    "1111111111100010",
    "1111111111100100",
    "1111111111100111",
    "1111111111101010",
    "1111111111101101",
    "1111111111110001",
    "1111111111110110",
    "1111111111111001",
    "1111111111111100",
    "1111111111111101",
    "1111111111111100",
    "1111111111111001",
    "1111111111110110",
    "1111111111110001",
    "1111111111101110",
    "1111111111101100",
    "1111111111101011",
    "1111111111101011",
    "1111111111101101",
    "1111111111101110",
    "1111111111110000",
    "1111111111110011",
    "1111111111110111",
    "1111111111111011",
    "1111111111111110",
    "1111111111111100",
    "1111111111111010",
    "1111111111111000",
    "1111111111110110",
    "1111111111110011",
    "1111111111101110",
    "1111111111101010",
    "1111111111100100",
    "1111111111100000",
    "1111111111011100",
    "1111111111011001",
    "1111111111010111",
    "1111111111011000",
    "1111111111011010",
    "1111111111011111",
    "1111111111100100",
    "1111111111101011",
    "1111111111110011",
    "1111111111111011",
    "1111111111111100",
    "1111111111110111",
    "1111111111110101",
    "1111111111110110",
    "1111111111111100",
    "1111111111111010",
    "1111111111110001",
    "1111111111101001",
    "1111111111100011",
    "1111111111100001",
    "1111111111100000",
    "1111111111100010",
    "1111111111100101",
    "1111111111101001",
    "1111111111101110",
    "1111111111110011",
    "1111111111111010",
    "1111111111111101",
    "1111111111111000",
    "1111111111110011",
    "1111111111110011",
    "1111111111110101",
    "1111111111111011",
    "1111111111111000",
    "1111111111101011",
    "1111111111011110",
    "1111111111001111",
    "1111111111000010",
    "1111111110110111",
    "1111111110110000",
    "1111111110101101",
    "1111111110101111",
    "1111111110110101",
    "1111111110111111",
    "1111111111001011",
    "1111111111011000",
    "1111111111100101",
    "1111111111110000",
    "1111111111111011",
    "1111111111111011",
    "1111111111110110",
    "1111111111110100",
    "1111111111110100",
    "1111111111111000",
    "1111111111111101",
    "1111111111111011",
    "1111111111110101",
    "1111111111110001",
    "1111111111101110",
    "1111111111101010",
    "1111111111100101",
    "1111111111011110",
    "1111111111010101",
    "1111111111010101",
    "1111111111101010",
    "1111111111011000",
    "1111111101101110",
    "1111111011011010",
    "1111111000101011",
    "1111110101111001",
    "1111110011011101",
    "1111110001100101",
    "1111110000011000",
    "1111101111110001",
    "1111101111101000",
    "1111101111111010",
    "1111110000100111",
    "1111110001110100",
    "1111110011100110",
    "1111110101111010",
    "1111111000101011",
    "1111111011101010",
    "1111111110100101",
    "1111111110110110",
    "1111111100111101",
    "1111111011110011",
    "1111111011001110",
    "1111111010111101",
    "1111111010101001",
    "1111111010000001",
    "1111111000111100",
    "1111110111011100",
    "1111110101101011",
    "1111110011111001",
    "1111110010010000",
    "1111110000110110",
    "1111101111101000",
    "1111101110011111",
    "1111101101011011",
    "1111101100100011",
    "1111101100000101",
    "1111101100010110",
    "1111101101100101",
    "1111101111110111",
    "1111110011000100",
    "1111110110110110",
    "1111111010110101",
    "1111111110101010",
    "1111111101110011",
    "1111111010110001",
    "1111111000001100",
    "1111110110000110",
    "1111110100011111",
    "1111110011011101",
    "1111110011000101",
    "1111110011100000",
    "1111110100110000",
    "1111110110101111",
    "1111111001001111",
    "1111111100000001",
    "1111111110110001",
    "1111111110101101",
    "1111111100100110",
    "1111111010110110",
    "1111111001010110",
    "1111110111111110",
    "1111110110100111",
    "1111110101010010",
    "1111110100000101",
    "1111110011001101",
    "1111110010110000",
    "1111110010110100",
    "1111110011001101",
    "1111110011101101",
    "1111110011111111",
    "1111110011111001",
    "1111110011011001",
    "1111110010101100",
    "1111110010001001",
    "1111110010000100",
    "1111110010101010",
    "1111110011111101",
    "1111110101110110",
    "1111111000000101",
    "1111111010011011",
    "1111111100110011",
    "1111111111001000",
    "1111111110011101",
    "1111111100000001",
    "1111111001100001",
    "1111110111000111",
    "1111110101000011",
    "1111110011100010",
    "1111110010110100",
    "1111110010111101",
    "1111110011111010",
    "1111110101100000",
    "1111110111100010",
    "1111111001110000",
    "1111111100000010",
    "1111111110010010",
    "1111111111011111",
    "1111111101011000",
    "1111111011010111",
    "1111111001100101",
    "1111111000001011",
    "1111110111010100",
    "1111110111000001",
    "1111110111001110",
    "1111110111110010",
    "1111111000011011",
    "1111111000111011",
    "1111111001001011",
    "1111111001001010",
    "1111111001000010",
    "1111111001000000",
    "1111111001001111",
    "1111111001110111",
    "1111111010110110",
    "1111111100000100",
    "1111111101011010",
    "1111111110110010",
    "1111111111110010",
    "1111111110010011",
    "1111111100101001",
    "1111111010110000",
    "1111111000101100",
    "1111110110100110",
    "1111110100101101",
    "1111110011010001",
    "1111110010011100",
    "1111110010010000",
    "1111110010101010",
    "1111110011011100",
    "1111110100011010",
    "1111110101011010",
    "1111110110010101",
    "1111110111001111",
    "1111111000001100",
    "1111111001001111",
    "1111111010011100",
    "1111111011110001",
    "1111111101001000",
    "1111111110011001",
    "1111111111100000",
    "1111111111100101",
    "1111111110111101",
    "1111111110100001",
    "1111111110001101",
    "1111111110000010",
    "1111111101111101",
    "1111111110000000",
    "1111111110001011",
    "1111111110100001",
    "1111111110111111",
    "1111111111100101",
    "1111111111101100",
    "1111111110111110",
    "1111111110001100",
    "1111111101011010",
    "1111111100101000",
    "1111111011111001",
    "1111111011001111",
    "1111111010101101",
    "1111111010010101",
    "1111111010000110",
    "1111111001111101",
    "1111111001111001",
    "1111111001110101",
    "1111111001101111",
    "1111111001100110",
    "1111111001011100",
    "1111111001010101",
    "1111111001011001",
    "1111111001101010",
    "1111111010001011",
    "1111111010111011",
    "1111111011110100",
    "1111111100101110",
    "1111111101100001",
    "1111111110000111",
    "1111111110011101",
    "1111111110101000",
    "1111111110101110",
    "1111111110111000",
    "1111111111001000",
    "1111111111011110",
    "1111111111110100",
    "1111111111111011",
    "1111111111111110",
    "1111111111100110",
    "1111111110111011",
    "1111111110000010",
    "1111111101000111",
    "1111111100010100",
    "1111111011101111",
    "1111111011011011",
    "1111111011010110",
    "1111111011011101",
    "1111111011100110",
    "1111111011101110",
    "1111111011101101",
    "1111111011100010",
    "1111111011001110",
    "1111111010110110",
    "1111111010100001",
    "1111111010011001",
    "1111111010100010",
    "1111111010111111",
    "1111111011101100",
    "1111111100011111",
    "1111111101001111",
    "1111111101110101",
    "1111111110001110",
    "1111111110011101",
    "1111111110101000",
    "1111111110110100",
    "1111111111001001",
    "1111111111100100",
    "1111111111111001",
    "1111111111011110",
    "1111111111001010",
    "1111111111000110",
    "1111111111010000",
    "1111111111100111",
    "1111111111111000",
    "1111111111011011",
    "1111111111000110",
    "1111111110111101",
    "1111111111000010",
    "1111111111010010",
    "1111111111101001",
    "1111111111111100",
    "1111111111101001",
    "1111111111100001",
    "1111111111100000",
    "1111111111100110",
    "1111111111101111",
    "1111111111110111",
    "1111111111111100",
    "1111111111111110",
    "1111111111111110",
    "1111111111111110",
    "1111111111111100",
    "1111111111111001",
    "1111111111110100",
    "1111111111110000",
    "1111111111101001",
    "1111111111100001",
    "1111111111010110",
    "1111111111000111",
    "1111111110110111",
    "1111111110101010",
    "1111111110100111",
    "1111111110110000",
    "1111111111001000",
    "1111111111101111",
    "1111111111011100",
    "1111111110100010",
    "1111111101101001",
    "1111111100110111",
    "1111111100010111",
    "1111111100001011",
    "1111111100010000",
    "1111111100100000",
    "1111111100101100",
    "1111111100101110",
    "1111111100100100",
    "1111111100010100",
    "1111111100000111",
    "1111111100001000",
    "1111111100011100",
    "1111111101000001",
    "1111111101110111",
    "1111111110110111",
    "1111111111111001",
    "1111111111000111",
    "1111111110010011",
    "1111111101101100",
    "1111111101010001",
    "1111111101000000",
    "1111111100110100",
    "1111111100101010",
    "1111111100011100",
    "1111111100001011",
    "1111111011111001",
    "1111111011101010",
    "1111111011100011",
    "1111111011100111",
    "1111111011111010",
    "1111111100011001",
    "1111111101000010",
    "1111111101101100",
    "1111111110001110",
    "1111111110100011",
    "1111111110100111",
    "1111111110011101",
    "1111111110001110",
    "1111111110000110",
    "1111111110001011",
    "1111111110100001",
    "1111111111000111",
    "1111111111110011",
    "1111111111100010",
    "1111111111000111",
    "1111111110111111",
    "1111111111001001",
    "1111111111011111",
    "1111111111111000",
    "1111111111101101",
    "1111111111011010",
    "1111111111001000",
    "1111111110110101",
    "1111111110011100",
    "1111111101111001",
    "1111111101001101",
    "1111111100011010",
    "1111111011100111",
    "1111111010111000",
    "1111111010010010",
    "1111111001110011",
    "1111111001011101",
    "1111111001001011",
    "1111111000111100",
    "1111111000110011",
    "1111111000110001",
    "1111111000111010",
    "1111111001010011",
    "1111111001111101",
    "1111111010111110",
    "1111111100010111",
    "1111111110001000",
    "1111111111110001",
    "1111111101100111",
    "1111111011100101",
    "1111111001111100",
    "1111111000111100",
    "1111111000101111",
    "1111111001011000",
    "1111111010110100",
    "1111111100110111",
    "1111111111010011",
    "1111111110000110",
    "1111111011100111",
    "1111111001011110",
    "1111110111110010",
    "1111110110100110",
    "1111110101111000",
    "1111110101100110",
    "1111110101100101",
    "1111110101101111",
    "1111110101111100",
    "1111110110000100",
    "1111110110000011",
    "1111110101110111",
    "1111110101100000",
    "1111110100111111",
    "1111110100011001",
    "1111110011110010",
    "1111110011010011",
    "1111110011000010",
    "1111110011001010",
    "1111110011110101",
    "1111110101000111",
    "1111110110111110",
    "1111111001010110",
    "1111111100000010",
    "1111111110110011",
    "1111111110100011",
    "1111111100010000",
    "1111111010011011",
    "1111111001000110",
    "1111111000010001",
    "1111110111110101",
    "1111110111101010",
    "1111110111101001",
    "1111110111101000",
    "1111110111100010",
    "1111110111010101",
    "1111110111000001",
    "1111110110101001",
    "1111110110010011",
    "1111110110000100",
    "1111110110000001",
    "1111110110001100",
    "1111110110100110",
    "1111110111010000",
    "1111111000001001",
    "1111111001001111",
    "1111111010011111",
    "1111111011110001",
    "1111111101000001",
    "1111111110000101",
    "1111111110111000",
    "1111111111010011",
    "1111111111010011",
    "1111111110111001",
    "1111111110000100",
    "1111111100111101",
    "1111111011101100",
    "1111111010100010",
    "1111111001101010",
    "1111111001010110",
    "1111111001101011",
    "1111111010101011",
    "1111111100001111",
    "1111111110001010",
    "1111111111110000",
    "1111111101110100",
    "1111111100001101",
    "1111111011000000",
    "1111111010010001",
    "1111111010000010",
    "1111111010010001",
    "1111111010111110",
    "1111111100000011",
    "1111111101011100",
    "1111111111000000",
    "1111111111011001",
    "1111111101111110",
    "1111111100110111",
    "1111111100001100",
    "1111111011111111",
    "1111111100001110",
    "1111111100110100",
    "1111111101100111",
    "1111111110011110",
    "1111111111010000",
    "1111111111111011",
    "1111111111100011",
    "1111111111001100",
    "1111111110111110",
    "1111111110110010",
    "1111111110101001",
    "1111111110100001",
    "1111111110011001",
    "1111111110010010",
    "1111111110001100",
    "1111111110001000",
    "1111111110000101",
    "1111111110000011",
    "1111111110000000",
    "1111111101111011",
    "1111111101110010",
    "1111111101100110",
    "1111111101010010",
    "1111111100110111",
    "1111111100010010",
    "1111111011011111",
    "1111111010100001",
    "1111111001010101",
    "1111111000000011",
    "1111110110110000",
    "1111110101100011",
    "1111110100100011",
    "1111110011111010",
    "1111110011101100",
    "1111110011111101",
    "1111110100110001",
    "1111110110000011",
    "1111110111110010",
    "1111111001110100",
    "1111111100000001",
    "1111111110001101",
    "1111111111101100",
    "1111111101111001",
    "1111111100011101",
    "1111111011011010",
    "1111111010110001",
    "1111111010100100",
    "1111111010110000",
    "1111111011010011",
    "1111111100000110",
    "1111111101000101",
    "1111111110001001",
    "1111111111001110",
    "1111111111101001",
    "1111111110100111",
    "1111111101100111",
    "1111111100101100",
    "1111111011111010",
    "1111111011010100",
    "1111111010111011",
    "1111111010101110",
    "1111111010101011",
    "1111111010101100",
    "1111111010101001",
    "1111111010011011",
    "1111111010000000",
    "1111111001010111",
    "1111111000100110",
    "1111110111110100",
    "1111110111001000",
    "1111110110101100",
    "1111110110100010",
    "1111110110101111",
    "1111110111010001",
    "1111111000001000",
    "1111111001010101",
    "1111111010110101",
    "1111111100100110",
    "1111111110100111",
    "1111111111001010",
    "1111111100111100",
    "1111111010110010",
    "1111111000110111",
    "1111110111010011",
    "1111110110001111",
    "1111110101101100",
    "1111110101101010",
    "1111110110000011",
    "1111110110110011",
    "1111110111110010",
    "1111111000111010",
    "1111111010000110",
    "1111111011010101",
    "1111111100100011",
    "1111111101101111",
    "1111111110110101",
    "1111111111110100",
    "1111111111010011",
    "1111111110101001",
    "1111111110000110",
    "1111111101101001",
    "1111111101001111",
    "1111111100110111",
    "1111111100100010",
    "1111111100010000",
    "1111111100000011",
    "1111111011111011",
    "1111111011111011",
    "1111111100000001",
    "1111111100001101",
    "1111111100011100",
    "1111111100101010",
    "1111111100111001",
    "1111111101001000",
    "1111111101011101",
    "1111111101111110",
    "1111111110101100",
    "1111111111101001",
    "1111111111001010",
    "1111111101111010",
    "1111111100100111",
    "1111111011010110",
    "1111111010001100",
    "1111111001001100",
    "1111111000011011",
    "1111110111111100",
    "1111110111101110",
    "1111110111110011",
    "1111111000000110",
    "1111111000101000",
    "1111111001010101",
    "1111111010001101",
    "1111111011001001",
    "1111111100000010",
    "1111111100110001",
    "1111111101010000",
    "1111111101011100",
    "1111111101011001",
    "1111111101001011",
    "1111111100111011",
    "1111111100110000",
    "1111111100101110",
    "1111111100111010",
    "1111111101010001",
    "1111111101110000",
    "1111111110010010",
    "1111111110110010",
    "1111111111001011",
    "1111111111011010",
    "1111111111011100",
    "1111111111010001",
    "1111111110111001",
    "1111111110010100",
    "1111111101100100",
    "1111111100101000",
    "1111111011100001",
    "1111111010010110",
    "1111111001001011",
    "1111111000001010",
    "1111110111011100",
    "1111110111001001",
    "1111110111010011",
    "1111110111111001",
    "1111111000110110",
    "1111111001111110",
    "1111111011000111",
    "1111111100000111",
    "1111111100110110",
    "1111111101010100",
    "1111111101100100",
    "1111111101101100",
    "1111111101110110",
    "1111111110001000",
    "1111111110100010",
    "1111111111000100",
    "1111111111100110",
    "1111111111111001",
    "1111111111100010",
    "1111111111010110",
    "1111111111010001",
    "1111111111010100",
    "1111111111011100",
    "1111111111100111",
    "1111111111111000",
    "1111111111101101",
    "1111111111001101",
    "1111111110100110",
    "1111111101111010",
    "1111111101010001",
    "1111111100110001",
    "1111111100011111",
    "1111111100011011",
    "1111111100100100",
    "1111111100110101",
    "1111111101001001",
    "1111111101011100",
    "1111111101110000",
    "1111111110001000",
    "1111111110100011",
    "1111111111000000",
    "1111111111011001",
    "1111111111101000",
    "1111111111101010",
    "1111111111011110",
    "1111111111001001",
    "1111111110110101",
    "1111111110101110",
    "1111111110111011",
    "1111111111011100",
    "1111111111110000",
    "1111111110111010",
    "1111111110001100",
    "1111111101101111",
    "1111111101101001",
    "1111111101111010",
    "1111111110100000",
    "1111111111010011",
    "1111111111101001",
    "1111111110011111",
    "1111111101001000",
    "1111111011100111",
    "1111111010000000",
    "1111111000011001",
    "1111110110111010",
    "1111110101101110",
    "1111110100111100",
    "1111110100101000",
    "1111110100110101",
    "1111110101100010",
    "1111110110101000",
    "1111110111111111",
    "1111111001011100",
    "1111111010110011",
    "1111111011111001",
    "1111111100101010",
    "1111111101000110",
    "1111111101010001",
    "1111111101010011",
    "1111111101011000",
    "1111111101100101",
    "1111111101111101",
    "1111111110100011",
    "1111111111010000",
    "1111111111111011",
    "1111111111000111",
    "1111111110011000",
    "1111111101101111",
    "1111111101001010",
    "1111111100101001",
    "1111111100001001",
    "1111111011101001",
    "1111111011001000",
    "1111111010101000",
    "1111111010001100",
    "1111111001111010",
    "1111111001110011",
    "1111111001111100",
    "1111111010001111",
    "1111111010101101",
    "1111111011010010",
    "1111111011111011",
    "1111111100100111",
    "1111111101010110",
    "1111111110000110",
    "1111111110110100",
    "1111111111011101",
    "1111111111111000",
    "1111111111111100",
    "1111111111110010",
    "1111111111001100",
    "1111111110010000",
    "1111111101000111",
    "1111111011111011",
    "1111111010111010",
    "1111111010010001",
    "1111111010001101",
    "1111111010110010",
    "1111111100000001",
    "1111111101110000",
    "1111111111110100",
    "1111111110000011",
    "1111111100001100",
    "1111111010110000",
    "1111111001111010",
    "1111111001101010",
    "1111111010000010",
    "1111111010111000",
    "1111111100000101",
    "1111111101011101",
    "1111111110110101",
    "1111111111111001",
    "1111111110111101",
    "1111111110010011",
    "1111111110000001",
    "1111111110000010",
    "1111111110010010",
    "1111111110101101",
    "1111111111001110",
    "1111111111101110",
    "1111111111110100",
    "1111111111100110",
    "1111111111101010",
    "1111111111110100",
    "1111111110111001",
    "1111111101011110",
    "1111111011101001",
    "1111111001100110",
    "1111110111100011",
    "1111110101110111",
    "1111110100110000",
    "1111110100011100",
    "1111110100111101",
    "1111110110010001",
    "1111111000001010",
    "1111111010010111",
    "1111111100100110",
    "1111111110101001",
    "1111111111100111",
    "1111111110010010",
    "1111111101010111",
    "1111111100101111",
    "1111111100011001",
    "1111111100010011",
    "1111111100011001",
    "1111111100101001",
    "1111111100111110",
    "1111111101010001",
    "1111111101011001",
    "1111111101001101",
    "1111111100101011",
    "1111111011110111",
    "1111111010110110",
    "1111111001110111",
    "1111111001000101",
    "1111111000101010",
    "1111111000101101",
    "1111111001001110",
    "1111111010001110",
    "1111111011100100",
    "1111111101001000",
    "1111111110101101",
    "1111111111110100",
    "1111111110110000",
    "1111111110001010",
    "1111111110000100",
    "1111111110011110",
    "1111111111010000",
    "1111111111101011",
    "1111111110101000",
    "1111111101101101",
    "1111111101000101",
    "1111111100110100",
    "1111111100111010",
    "1111111101010011",
    "1111111101111001",
    "1111111110100111",
    "1111111111010101",
    "1111111111111011",
    "1111111111010001",
    "1111111110101100",
    "1111111110001111",
    "1111111101111101",
    "1111111101111100",
    "1111111110010001",
    "1111111110111101",
    "1111111111111100",
    "1111111110110110",
    "1111111101101011",
    "1111111100101010",
    "1111111011111110",
    "1111111011101101",
    "1111111011110111",
    "1111111100011010",
    "1111111101001111",
    "1111111110001101",
    "1111111111001101",
    "1111111111110011",
    "1111111110111010",
    "1111111110000101",
    "1111111101010010",
    "1111111100100011",
    "1111111011111010",
    "1111111011011100",
    "1111111011001101",
    "1111111011010011",
    "1111111011101101",
    "1111111100011010",
    "1111111101010110",
    "1111111110010111",
    "1111111111010100",
    "1111111111111100",
    "1111111111100111",
    "1111111111101110",
    "1111111111101101",
    "1111111110110101",
    "1111111101110000",
    "1111111100100110",
    "1111111011011101",
    "1111111010011101",
    "1111111001101010",
    "1111111001000100",
    "1111111000101011",
    "1111111000011011",
    "1111111000010000",
    "1111111000001000",
    "1111111000000000",
    "1111110111111101",
    "1111110111111101",
    "1111111000000010",
    "1111111000001011",
    "1111111000010101",
    "1111111000011101",
    "1111111000100001",
    "1111111000011111",
    "1111111000011001",
    "1111111000010010",
    "1111111000010000",
    "1111111000010011",
    "1111111000100011",
    "1111111000111110",
    "1111111001100100",
    "1111111010010010",
    "1111111011000011",
    "1111111011110011",
    "1111111100100000",
    "1111111101000111",
    "1111111101101011",
    "1111111110001101",
    "1111111110101111",
    "1111111111001111",
    "1111111111101101",
    "1111111111111000",
    "1111111111101001",
    "1111111111100100",
    "1111111111101101",
    "1111111111111001",
    "1111111111010010",
    "1111111110011001",
    "1111111101001111",
    "1111111011110111",
    "1111111010010110",
    "1111111000110110",
    "1111110111011111",
    "1111110110011010",
    "1111110101101011",
    "1111110101010010",
    "1111110101001110",
    "1111110101011001",
    "1111110101110000",
    "1111110110010000",
    "1111110110110111",
    "1111110111101000",
    "1111111000100101",
    "1111111001110000",
    "1111111011000100",
    "1111111100011110",
    "1111111101110011",
    "1111111110111100",
    "1111111111110011",
    "1111111111100110",
    "1111111111010011",
    "1111111111001100",
    "1111111111001100",
    "1111111111001111",
    "1111111111010011",
    "1111111111011001",
    "1111111111100001",
    "1111111111101111",
    "1111111111111011",
    "1111111111100010",
    "1111111111001010",
    "1111111110111001",
    "1111111110110011",
    "1111111110111100",
    "1111111111010001",
    "1111111111101101",
    "1111111111110110",
    "1111111111101001",
    "1111111111101100",
    "1111111111111000",
    "1111111111001101",
    "1111111110010110",
    "1111111101011100",
    "1111111100101001",
    "1111111100000101",
    "1111111011110110",
    "1111111011111011",
    "1111111100010100",
    "1111111100111010",
    "1111111101101010",
    "1111111110100001",
    "1111111111100000",
    "1111111111010101",
    "1111111110000100",
    "1111111100101101",
    "1111111011011001",
    "1111111010001111",
    "1111111001011000",
    "1111111000111001",
    "1111111000110010",
    "1111111001000000",
    "1111111001011001",
    "1111111001111000",
    "1111111010010010",
    "1111111010100110",
    "1111111010110010",
    "1111111010110110",
    "1111111010110110",
    "1111111010110101",
    "1111111010110100",
    "1111111010110110",
    "1111111011000000",
    "1111111011010011",
    "1111111011110100",
    "1111111100100110",
    "1111111101100101",
    "1111111110101111",
    "1111111111111010",
    "1111111110111111",
    "1111111110001011",
    "1111111101101011",
    "1111111101100011",
    "1111111101101110",
    "1111111110001000",
    "1111111110101011",
    "1111111111010010",
    "1111111111111000",
    "1111111111100010",
    "1111111111000010",
    "1111111110100010",
    "1111111110000011",
    "1111111101100001",
    "1111111100111101",
    "1111111100011001",
    "1111111011110101",
    "1111111011010100",
    "1111111010110110",
    "1111111010011001",
    "1111111001111100",
    "1111111001011110",
    "1111111000111100",
    "1111111000011100",
    "1111111000000000",
    "1111110111110000",
    "1111110111101111",
    "1111111000000001",
    "1111111000100111",
    "1111111001011101",
    "1111111010011100",
    "1111111011100000",
    "1111111100100100",
    "1111111101100011",
    "1111111110011011",
    "1111111111001010",
    "1111111111110010",
    "1111111111101010",
    "1111111111001110",
    "1111111110110111",
    "1111111110100011",
    "1111111110010001",
    "1111111110000101",
    "1111111101111101",
    "1111111101111001",
    "1111111101110111",
    "1111111101110100",
    "1111111101101111",
    "1111111101101000",
    "1111111101100011",
    "1111111101100110",
    "1111111101111000",
    "1111111110011111",
    "1111111111011101",
    "1111111111001001",
    "1111111101011111",
    "1111111011100111",
    "1111111001101101",
    "1111110111111011",
    "1111110110011011",
    "1111110101010011",
    "1111110100101001",
    "1111110100011110",
    "1111110100110000",
    "1111110101011011",
    "1111110110011001",
    "1111110111100100",
    "1111111000110110",
    "1111111010001000",
    "1111111011010011",
    "1111111100010001",
    "1111111100111100",
    "1111111101010001",
    "1111111101010000",
    "1111111100111101",
    "1111111100011110",
    "1111111011111011",
    "1111111011011110",
    "1111111011001101",
    "1111111011001011",
    "1111111011011001",
    "1111111011110100",
    "1111111100011101",
    "1111111101001111",
    "1111111110001000",
    "1111111111000110",
    "1111111111110101",
    "1111111110110101",
    "1111111101111100",
    "1111111101001111",
    "1111111100110011",
    "1111111100101100",
    "1111111100111101",
    "1111111101100101",
    "1111111110100100",
    "1111111111110111",
    "1111111110100011",
    "1111111100110110",
    "1111111011001000",
    "1111111001011111",
    "1111111000000100",
    "1111110110111111",
    "1111110110010101",
    "1111110110001011",
    "1111110110100100",
    "1111110111011011",
    "1111111000101101",
    "1111111010001110",
    "1111111011110001",
    "1111111101001101",
    "1111111110010110",
    "1111111111000111",
    "1111111111011110",
    "1111111111011100",
    "1111111111001001",
    "1111111110101100",
    "1111111110001101",
    "1111111101110010",
    "1111111101100001",
    "1111111101100000",
    "1111111101110010",
    "1111111110011001",
    "1111111111010111",
    "1111111111010101",
    "1111111101110100",
    "1111111100001101",
    "1111111010101001",
    "1111111001010011",
    "1111111000010011",
    "1111110111110010",
    "1111110111110001",
    "1111111000001110",
    "1111111001000101",
    "1111111010010000",
    "1111111011100110",
    "1111111100111110",
    "1111111110010101",
    "1111111111100010",
    "1111111111011101",
    "1111111110110010",
    "1111111110100000",
    "1111111110100101",
    "1111111111000000",
    "1111111111101001",
    "1111111111100010",
    "1111111110110000",
    "1111111110000111",
    "1111111101101100",
    "1111111101100100",
    "1111111101101111",
    "1111111110001001",
    "1111111110101101",
    "1111111111010010",
    "1111111111110001",
    "1111111111111000",
    "1111111111110110",
    "1111111111111000",
    "1111111111010101",
    "1111111110100010",
    "1111111101100110",
    "1111111100100110",
    "1111111011101010",
    "1111111010111000",
    "1111111010010110",
    "1111111010000101",
    "1111111010000101",
    "1111111010010110",
    "1111111010110011",
    "1111111011011001",
    "1111111100000011",
    "1111111100101101",
    "1111111101010011",
    "1111111101110001",
    "1111111110000111",
    "1111111110010110",
    "1111111110100001",
    "1111111110101010",
    "1111111110110111",
    "1111111111001100",
    "1111111111101101",
    "1111111111100010",
    "1111111110101011",
    "1111111101101101",
    "1111111100101101",
    "1111111011110100",
    "1111111011001000",
    "1111111010101100",
    "1111111010100011",
    "1111111010101101",
    "1111111011001001",
    "1111111011110010",
    "1111111100100011",
    "1111111101011000",
    "1111111110001010",
    "1111111110110111",
    "1111111111011100",
    "1111111111110111",
    "1111111111110100",
    "1111111111101001",
    "1111111111100101",
    "1111111111100011",
    "1111111111100100",
    "1111111111100110",
    "1111111111101001",
    "1111111111101100",
    "1111111111110000",
    "1111111111110000",
    "1111111111101010",
    "1111111111011111",
    "1111111111001001",
    "1111111110101011",
    "1111111110000110",
    "1111111101011110",
    "1111111100111001",
    "1111111100011010",
    "1111111100000110",
    "1111111100000001",
    "1111111100001010",
    "1111111100100010",
    "1111111101001001",
    "1111111101111100",
    "1111111110111001",
    "1111111111111011",
    "1111111110111101",
    "1111111101111001",
    "1111111100111011",
    "1111111100000111",
    "1111111011100011",
    "1111111011010001",
    "1111111011010101",
    "1111111011101111",
    "1111111100011000",
    "1111111101001011",
    "1111111101111110",
    "1111111110101001",
    "1111111111000101",
    "1111111111010000",
    "1111111111001100",
    "1111111110111110",
    "1111111110101001",
    "1111111110010000",
    "1111111101111000",
    "1111111101100100",
    "1111111101010010",
    "1111111101000111",
    "1111111101000100",
    "1111111101001011",
    "1111111101011110",
    "1111111101111110",
    "1111111110101011",
    "1111111111100011",
    "1111111111011101",
    "1111111110011110",
    "1111111101100011",
    "1111111100110001",
    "1111111100001001",
    "1111111011110000",
    "1111111011100110",
    "1111111011101101",
    "1111111100000011",
    "1111111100100100",
    "1111111101001111",
    "1111111101111101",
    "1111111110101001",
    "1111111111001111",
    "1111111111101000",
    "1111111111110100",
    "1111111111110001",
    "1111111111100000",
    "1111111111000011",
    "1111111110011111",
    "1111111101110111",
    "1111111101010000",
    "1111111100101100",
    "1111111100001111",
    "1111111011111100",
    "1111111011110101",
    "1111111011111010",
    "1111111100001101",
    "1111111100101100",
    "1111111101011001",
    "1111111110010000",
    "1111111111001111",
    "1111111111101100",
    "1111111110101111",
    "1111111101111111",
    "1111111101100011",
    "1111111101011110",
    "1111111101110011",
    "1111111110100001",
    "1111111111011111",
    "1111111111010110",
    "1111111110001001",
    "1111111100111101",
    "1111111011110011",
    "1111111010101100",
    "1111111001101001",
    "1111111000101100",
    "1111110111111000",
    "1111110111010101",
    "1111110111000101",
    "1111110111001101",
    "1111110111101010",
    "1111111000011000",
    "1111111001001100",
    "1111111001111100",
    "1111111010100010",
    "1111111010110110",
    "1111111010111101",
    "1111111010111000",
    "1111111010101111",
    "1111111010101010",
    "1111111010101100",
    "1111111010111011",
    "1111111011010100",
    "1111111011110111",
    "1111111100100000",
    "1111111101001010",
    "1111111101110100",
    "1111111110011110",
    "1111111111000111",
    "1111111111101111",
    "1111111111100110",
    "1111111111000001",
    "1111111110100001",
    "1111111110001001",
    "1111111101111011",
    "1111111101111011",
    "1111111110001001",
    "1111111110100001",
    "1111111111000011",
    "1111111111101101",
    "1111111111011101",
    "1111111110100010",
    "1111111101011111",
    "1111111100010110",
    "1111111011001010",
    "1111111010000010",
    "1111111001000010",
    "1111111000001111",
    "1111110111101100",
    "1111110111011101",
    "1111110111011111",
    "1111110111110000",
    "1111111000001110",
    "1111111000110100",
    "1111111001100010",
    "1111111010010111",
    "1111111011010001",
    "1111111100001111",
    "1111111101010010",
    "1111111110010111",
    "1111111111011011",
    "1111111111100010",
    "1111111110100101",
    "1111111101101101",
    "1111111100110111",
    "1111111100000101",
    "1111111011010101",
    "1111111010101010",
    "1111111010000011",
    "1111111001100101",
    "1111111001010010",
    "1111111001001111",
    "1111111001011100",
    "1111111001111001",
    "1111111010100011",
    "1111111011010100",
    "1111111100001100",
    "1111111101000101",
    "1111111110000000",
    "1111111110111101",
    "1111111111111100",
    "1111111111000000",
    "1111111101111110",
    "1111111100111111",
    "1111111100001001",
    "1111111011011111",
    "1111111011000111",
    "1111111010111110",
    "1111111011000110",
    "1111111011011000",
    "1111111011110001",
    "1111111100001101",
    "1111111100100110",
    "1111111100111100",
    "1111111101001110",
    "1111111101011101",
    "1111111101101110",
    "1111111110000011",
    "1111111110011111",
    "1111111111000011",
    "1111111111101111",
    "1111111111011101",
    "1111111110101000",
    "1111111101110011",
    "1111111101000000",
    "1111111100010000",
    "1111111011100100",
    "1111111010111111",
    "1111111010100001",
    "1111111010001101",
    "1111111010000011",
    "1111111010000100",
    "1111111010001111",
    "1111111010100011",
    "1111111010111111",
    "1111111011011111",
    "1111111100000011",
    "1111111100101010",
    "1111111101010010",
    "1111111101111101",
    "1111111110101010",
    "1111111111011011",
    "1111111111101110",
    "1111111110111001",
    "1111111110000100",
    "1111111101010011",
    "1111111100101010",
    "1111111100001101",
    "1111111100000000",
    "1111111100000110",
    "1111111100100001",
    "1111111101001110",
    "1111111110001001",
    "1111111111001101",
    "1111111111100111",
    "1111111110011110",
    "1111111101010111",
    "1111111100010110",
    "1111111011011101",
    "1111111010101110",
    "1111111010001100",
    "1111111001110100",
    "1111111001100110",
    "1111111001011110",
    "1111111001011001",
    "1111111001010111",
    "1111111001011000",
    "1111111001011110",
    "1111111001101001",
    "1111111001111100",
    "1111111010010011",
    "1111111010101101",
    "1111111011000110",
    "1111111011011001",
    "1111111011100100",
    "1111111011101000",
    "1111111011101010",
    "1111111011101101",
    "1111111011110110",
    "1111111100001010",
    "1111111100101011",
    "1111111101011010",
    "1111111110010011",
    "1111111111010011",
    "1111111111101010",
    "1111111110101111",
    "1111111101111110",
    "1111111101010111",
    "1111111100111011",
    "1111111100101010",
    "1111111100100100",
    "1111111100101010",
    "1111111100111001",
    "1111111101010100",
    "1111111101111000",
    "1111111110100101",
    "1111111111010101",
    "1111111111110110",
    "1111111111001000",
    "1111111110011110",
    "1111111101111001",
    "1111111101011000",
    "1111111100111001",
    "1111111100011010",
    "1111111011111101",
    "1111111011100001",
    "1111111011001000",
    "1111111010110011",
    "1111111010100011",
    "1111111010011001",
    "1111111010010011",
    "1111111010010011",
    "1111111010010110",
    "1111111010011010",
    "1111111010100000",
    "1111111010100111",
    "1111111010110001",
    "1111111010111110",
    "1111111011001101",
    "1111111011100000",
    "1111111011110101",
    "1111111100001001",
    "1111111100010111",
    "1111111100100000",
    "1111111100100010",
    "1111111100011101",
    "1111111100010001",
    "1111111100000001",
    "1111111011101100",
    "1111111011010100",
    "1111111010111110",
    "1111111010101001",
    "1111111010011011",
    "1111111010010110",
    "1111111010011011",
    "1111111010101010",
    "1111111011000001",
    "1111111011011111",
    "1111111100000000",
    "1111111100100011",
    "1111111101001001",
    "1111111101110100",
    "1111111110100100",
    "1111111111011011",
    "1111111111100111",
    "1111111110101101",
    "1111111101111000",
    "1111111101010001",
    "1111111100111110",
    "1111111101000001",
    "1111111101011101",
    "1111111110001101",
    "1111111111001100",
    "1111111111101001",
    "1111111110100001",
    "1111111101100000",
    "1111111100101110",
    "1111111100001111",
    "1111111100000100",
    "1111111100001101",
    "1111111100100111",
    "1111111101001100",
    "1111111101111000",
    "1111111110101000",
    "1111111111011001",
    "1111111111110010",
    "1111111110111110",
    "1111111110000111",
    "1111111101001110",
    "1111111100010111",
    "1111111011100011",
    "1111111010110110",
    "1111111010010100",
    "1111111001111101",
    "1111111001110010",
    "1111111001110011",
    "1111111010000001",
    "1111111010011010",
    "1111111010111110",
    "1111111011101010",
    "1111111100011101",
    "1111111101010000",
    "1111111101111111",
    "1111111110100111",
    "1111111111000100",
    "1111111111010110",
    "1111111111011110",
    "1111111111011111",
    "1111111111011101",
    "1111111111011011",
    "1111111111011010",
    "1111111111011010",
    "1111111111011011",
    "1111111111011010",
    "1111111111011001",
    "1111111111010111",
    "1111111111010101",
    "1111111111010100",
    "1111111111010011",
    "1111111111010010",
    "1111111111001111",
    "1111111111000110",
    "1111111110110110",
    "1111111110100001",
    "1111111110000110",
    "1111111101101001",
    "1111111101001110",
    "1111111100110111",
    "1111111100100110",
    "1111111100011000",
    "1111111100001110",
    "1111111100000011",
    "1111111011110110",
    "1111111011100101",
    "1111111011010011",
    "1111111011000010",
    "1111111010110110",
    "1111111010101111",
    "1111111010101111",
    "1111111010110101",
    "1111111011000000",
    "1111111011001011",
    "1111111011010101",
    "1111111011011101",
    "1111111011100011",
    "1111111011101001",
    "1111111011110011",
    "1111111100000010",
    "1111111100010111",
    "1111111100110010",
    "1111111101010001",
    "1111111101110000",
    "1111111110001101",
    "1111111110101001",
    "1111111111000011",
    "1111111111011100",
    "1111111111110110",
    "1111111111101101",
    "1111111111010011",
    "1111111110111011",
    "1111111110100110",
    "1111111110010110",
    "1111111110001100",
    "1111111110000110",
    "1111111110000011",
    "1111111110000010",
    "1111111110000101",
    "1111111110001010",
    "1111111110010011",
    "1111111110100011",
    "1111111110111000",
    "1111111111010010",
    "1111111111110011",
    "1111111111101001",
    "1111111111001000",
    "1111111110101100",
    "1111111110010101",
    "1111111110000110",
    "1111111101111101",
    "1111111101111000",
    "1111111101110111",
    "1111111101110110",
    "1111111101110101",
    "1111111101110101",
    "1111111101110111",
    "1111111101111010",
    "1111111110000000",
    "1111111110000110",
    "1111111110001011",
    "1111111110001011",
    "1111111110000011",
    "1111111101110011",
    "1111111101011100",
    "1111111101000010",
    "1111111100101001",
    "1111111100010101",
    "1111111100001010",
    "1111111100001011",
    "1111111100011001",
    "1111111100110101",
    "1111111101011101",
    "1111111110010000",
    "1111111111001100",
    "1111111111101101",
    "1111111110100111",
    "1111111101100001",
    "1111111100011111",
    "1111111011100111",
    "1111111011000000",
    "1111111010101111",
    "1111111010111000",
    "1111111011011100",
    "1111111100011000",
    "1111111101100110",
    "1111111110111101",
    "1111111111101001",
    "1111111110011100",
    "1111111101011100",
    "1111111100101101",
    "1111111100001110",
    "1111111100000000",
    "1111111100000001",
    "1111111100001111",
    "1111111100101100",
    "1111111101010100",
    "1111111110000100",
    "1111111110111000",
    "1111111111101000",
    "1111111111101011",
    "1111111111001101",
    "1111111110111100",
    "1111111110110110",
    "1111111110111000",
    "1111111111000000",
    "1111111111001001",
    "1111111111010001",
    "1111111111010110",
    "1111111111010101",
    "1111111111001110",
    "1111111110111111",
    "1111111110100111",
    "1111111110001000",
    "1111111101100100",
    "1111111100111101",
    "1111111100011001",
    "1111111011111010",
    "1111111011100000",
    "1111111011001100",
    "1111111011000000",
    "1111111010111101",
    "1111111011000010",
    "1111111011010011",
    "1111111011110000",
    "1111111100010111",
    "1111111101001011",
    "1111111110001000",
    "1111111111001011",
    "1111111111101001",
    "1111111110100000",
    "1111111101011001",
    "1111111100011011",
    "1111111011101001",
    "1111111011000110",
    "1111111010110000",
    "1111111010100110",
    "1111111010100011",
    "1111111010100011",
    "1111111010100000",
    "1111111010011001",
    "1111111010001101",
    "1111111001111110",
    "1111111001101101",
    "1111111001011110",
    "1111111001001111",
    "1111111001000011",
    "1111111000111010",
    "1111111000110101",
    "1111111000110011",
    "1111111000110110",
    "1111111001000001",
    "1111111001011000",
    "1111111001111110",
    "1111111010110110",
    "1111111011111110",
    "1111111101010101",
    "1111111110110101",
    "1111111111100011",
    "1111111110000001",
    "1111111100100110",
    "1111111011010111",
    "1111111010011000",
    "1111111001101101",
    "1111111001011000",
    "1111111001011010",
    "1111111001110011",
    "1111111010100000",
    "1111111011011110",
    "1111111100101010",
    "1111111101111101",
    "1111111111010010",
    "1111111111010111",
    "1111111110001011",
    "1111111101001001",
    "1111111100011000",
    "1111111011111000",
    "1111111011101011",
    "1111111011110001",
    "1111111100001000",
    "1111111100101011",
    "1111111101010111",
    "1111111110000101",
    "1111111110101111",
    "1111111111010101",
    "1111111111110100",
    "1111111111101110",
    "1111111111011001",
    "1111111111000101",
    "1111111110110011",
    "1111111110100011",
    "1111111110010001",
    "1111111101111101",
    "1111111101100110",
    "1111111101001001",
    "1111111100100110",
    "1111111011111010",
    "1111111011000110",
    "1111111010001001",
    "1111111001000101",
    "1111110111111111",
    "1111110110111011",
    "1111110110000001",
    "1111110101011000",
    "1111110101000100",
    "1111110101001101",
    "1111110101110011",
    "1111110110110101",
    "1111111000001111",
    "1111111001111010",
    "1111111011101100",
    "1111111101011100",
    "1111111111000011",
    "1111111111100100",
    "1111111110011111",
    "1111111101101101",
    "1111111101001101",
    "1111111100111110",
    "1111111100111111",
    "1111111101010000",
    "1111111101101110",
    "1111111110010101",
    "1111111111000000",
    "1111111111100111",
    "1111111111111000",
    "1111111111100110",
    "1111111111100010",
    "1111111111100101",
    "1111111111101011",
    "1111111111101110",
    "1111111111101001",
    "1111111111011011",
    "1111111111000100",
    "1111111110100110",
    "1111111110000110",
    "1111111101100111",
    "1111111101001001",
    "1111111100110001",
    "1111111100011101",
    "1111111100001101",
    "1111111100000001",
    "1111111011111001",
    "1111111011110110",
    "1111111011111001",
    "1111111100000010",
    "1111111100010101",
    "1111111100110001",
    "1111111101011000",
    "1111111110000111",
    "1111111110111100",
    "1111111111110110",
    "1111111111001101",
    "1111111110010100",
    "1111111101011110",
    "1111111100110000",
    "1111111100001011",
    "1111111011110011",
    "1111111011101010",
    "1111111011110001",
    "1111111100000111",
    "1111111100101001",
    "1111111101010010",
    "1111111101111110",
    "1111111110101100",
    "1111111111011010",
    "1111111111110110",
    "1111111111000111",
    "1111111110011000",
    "1111111101101001",
    "1111111100111010",
    "1111111100010000",
    "1111111011101101",
    "1111111011010011",
    "1111111011000010",
    "1111111010111000",
    "1111111010110010",
    "1111111010101100",
    "1111111010100100",
    "1111111010011100",
    "1111111010010110",
    "1111111010010010",
    "1111111010010100",
    "1111111010011101",
    "1111111010101100",
    "1111111011000000",
    "1111111011010110",
    "1111111011110010",
    "1111111100010010",
    "1111111100111000",
    "1111111101100100",
    "1111111110010101",
    "1111111111001001",
    "1111111111111101",
    "1111111111010000",
    "1111111110101000",
    "1111111110001000",
    "1111111101110001",
    "1111111101100110",
    "1111111101100111",
    "1111111101110011",
    "1111111110001100",
    "1111111110101101",
    "1111111111010111",
    "1111111111111000",
    "1111111111000101",
    "1111111110001111",
    "1111111101010111",
    "1111111100100000",
    "1111111011101010",
    "1111111010111010",
    "1111111010010101",
    "1111111001111100",
    "1111111001110100",
    "1111111001111100",
    "1111111010010101",
    "1111111010111100",
    "1111111011101110",
    "1111111100100110",
    "1111111101011101",
    "1111111110010000",
    "1111111110111011",
    "1111111111011101",
    "1111111111111001",
    "1111111111101000",
    "1111111111001101",
    "1111111110101110",
    "1111111110001101",
    "1111111101101010",
    "1111111101000110",
    "1111111100100000",
    "1111111011110110",
    "1111111011000111",
    "1111111010010010",
    "1111111001011000",
    "1111111000011110",
    "1111110111101001",
    "1111110110111110",
    "1111110110100011",
    "1111110110011001",
    "1111110110100000",
    "1111110110110111",
    "1111110111011010",
    "1111111000001001",
    "1111111001000010",
    "1111111010000011",
    "1111111011001011",
    "1111111100010111",
    "1111111101100000",
    "1111111110100001",
    "1111111111010010",
    "1111111111101110",
    "1111111111110110",
    "1111111111101001",
    "1111111111001101",
    "1111111110101000",
    "1111111101111100",
    "1111111101001110",
    "1111111100011110",
    "1111111011101110",
    "1111111010111111",
    "1111111010010100",
    "1111111001110000",
    "1111111001010101",
    "1111111001000111",
    "1111111001000101",
    "1111111001001111",
    "1111111001100001",
    "1111111001111000",
    "1111111010010000",
    "1111111010100111",
    "1111111010111100",
    "1111111011001111",
    "1111111011100011",
    "1111111011111000",
    "1111111100001111",
    "1111111100101010",
    "1111111101000111",
    "1111111101100111",
    "1111111110001000",
    "1111111110101001",
    "1111111111001010",
    "1111111111101100",
    "1111111111110001",
    "1111111111010011",
    "1111111110111000",
    "1111111110100001",
    "1111111110001101",
    "1111111101111111",
    "1111111101110111",
    "1111111101110101",
    "1111111101111010",
    "1111111110000101",
    "1111111110010100",
    "1111111110100110",
    "1111111110111011",
    "1111111111001110",
    "1111111111100001",
    "1111111111110000",
    "1111111111111100",
    "1111111111111011",
    "1111111111111011",
    "1111111111111100",
    "1111111111110000",
    "1111111111100000",
    "1111111111001100",
    "1111111110111001",
    "1111111110101001",
    "1111111110011110",
    "1111111110011000",
    "1111111110011001",
    "1111111110100000",
    "1111111110101010",
    "1111111110111000",
    "1111111111001001",
    "1111111111100001",
    "1111111111111110",
    "1111111111010111",
    "1111111110100100",
    "1111111101100110",
    "1111111100100001",
    "1111111011011010",
    "1111111010010110",
    "1111111001011110",
    "1111111000110100",
    "1111111000011011",
    "1111111000010010",
    "1111111000010100",
    "1111111000011011",
    "1111111000100011",
    "1111111000101001",
    "1111111000101100",
    "1111111000101101",
    "1111111000101110",
    "1111111000110011",
    "1111111000111111",
    "1111111001010100",
    "1111111001110001",
    "1111111010011001",
    "1111111011001100",
    "1111111100001001",
    "1111111101010000",
    "1111111110100000",
    "1111111111110110",
    "1111111110101010",
    "1111111101001011",
    "1111111011101011",
    "1111111010001101",
    "1111111000110101",
    "1111110111100111",
    "1111110110101000",
    "1111110101111010",
    "1111110101100100",
    "1111110101100100",
    "1111110101111101",
    "1111110110101011",
    "1111110111101110",
    "1111111001000000",
    "1111111010011001",
    "1111111011110000",
    "1111111100111101",
    "1111111101111001",
    "1111111110011111",
    "1111111110101101",
    "1111111110100101",
    "1111111110001010",
    "1111111101100001",
    "1111111100110000",
    "1111111011111001",
    "1111111010111111",
    "1111111010000011",
    "1111111001000111",
    "1111111000001110",
    "1111110111011100",
    "1111110110110100",
    "1111110110011010",
    "1111110110001011",
    "1111110110000111",
    "1111110110001011",
    "1111110110010010",
    "1111110110011010",
    "1111110110100010",
    "1111110110101010",
    "1111110110110001",
    "1111110110110111",
    "1111110110111000",
    "1111110110110001",
    "1111110110011111",
    "1111110110000101",
    "1111110101100100",
    "1111110101000001",
    "1111110100100111",
    "1111110100011010",
    "1111110100100001",
    "1111110100111111",
    "1111110101110100",
    "1111110110111011",
    "1111111000010100",
    "1111111001111000",
    "1111111011100001",
    "1111111101001100",
    "1111111110110010",
    "1111111111101011",
    "1111111110010110",
    "1111111101001110",
    "1111111100010100",
    "1111111011101001",
    "1111111011001100",
    "1111111010111010",
    "1111111010101101",
    "1111111010100010",
    "1111111010010110",
    "1111111010001001",
    "1111111001111101",
    "1111111001111001",
    "1111111001111101",
    "1111111010010001",
    "1111111010110110",
    "1111111011101011",
    "1111111100101101",
    "1111111101110110",
    "1111111110111111",
    "1111111111111101",
    "1111111111001001",
    "1111111110100100",
    "1111111110001101",
    "1111111110000011",
    "1111111110000000",
    "1111111110000010",
    "1111111110000100",
    "1111111110000001",
    "1111111101111000",
    "1111111101100101",
    "1111111101000111",
    "1111111100011111",
    "1111111011101111",
    "1111111011000000",
    "1111111010011001",
    "1111111010000110",
    "1111111010001100",
    "1111111010110000",
    "1111111011110000",
    "1111111101000111",
    "1111111110101011",
    "1111111111100110",
    "1111111101111011",
    "1111111100010110",
    "1111111010111100",
    "1111111001101111",
    "1111111000110001",
    "1111111000000110",
    "1111110111101100",
    "1111110111100011",
    "1111110111101011",
    "1111111000000000",
    "1111111000100010",
    "1111111001001100",
    "1111111001111101",
    "1111111010110011",
    "1111111011101010",
    "1111111100100000",
    "1111111101010000",
    "1111111101111001",
    "1111111110011010",
    "1111111110110010",
    "1111111111000111",
    "1111111111011100",
    "1111111111110110",
    "1111111111100101",
    "1111111110111011",
    "1111111110001001",
    "1111111101010110",
    "1111111100100101",
    "1111111011111011",
    "1111111011011010",
    "1111111011000001",
    "1111111010110001",
    "1111111010101001",
    "1111111010100111",
    "1111111010110000",
    "1111111011000110",
    "1111111011101010",
    "1111111100100000",
    "1111111101100101",
    "1111111110110110",
    "1111111111101110",
    "1111111110010001",
    "1111111100110100",
    "1111111011011010",
    "1111111010001010",
    "1111111001001100",
    "1111111000100111",
    "1111111000011101",
    "1111111000110000",
    "1111111001011100",
    "1111111010010101",
    "1111111011010000",
    "1111111011111100",
    "1111111100010000",
    "1111111100000011",
    "1111111011010111",
    "1111111010001111",
    "1111111000111000",
    "1111110111011101",
    "1111110110001001",
    "1111110101000100",
    "1111110100010010",
    "1111110011110110",
    "1111110011101111",
    "1111110011111101",
    "1111110100100000",
    "1111110101010111",
    "1111110110011111",
    "1111110111110110",
    "1111111001010011",
    "1111111010101101",
    "1111111011111101",
    "1111111100111001",
    "1111111101011100",
    "1111111101100101",
    "1111111101010011",
    "1111111100101101",
    "1111111011111010",
    "1111111010111111",
    "1111111010000111",
    "1111111001010111",
    "1111111000110010",
    "1111111000011011",
    "1111111000010001",
    "1111111000010000",
    "1111111000010111",
    "1111111000100100",
    "1111111000110101",
    "1111111001000110",
    "1111111001011001",
    "1111111001101010",
    "1111111001111000",
    "1111111001111100",
    "1111111001110011",
    "1111111001011011",
    "1111111000110011",
    "1111111000000000",
    "1111110111001000",
    "1111110110010100",
    "1111110101101100",
    "1111110101011000",
    "1111110101011010",
    "1111110101110100",
    "1111110110101000",
    "1111110111110111",
    "1111111001100001",
    "1111111011100111",
    "1111111110000110",
    "1111111111000011",
    "1111111100000001",
    "1111111000111001",
    "1111110101110110",
    "1111110011000010",
    "1111110000101011",
    "1111101110111010",
    "1111101101110111",
    "1111101101100101",
    "1111101110000011",
    "1111101111001011",
    "1111110000110001",
    "1111110010101110",
    "1111110100111010",
    "1111110111001110",
    "1111111001100001",
    "1111111011101110",
    "1111111101101100",
    "1111111111010101",
    "1111111111010111",
    "1111111110011011",
    "1111111101110000",
    "1111111101001110",
    "1111111100101111",
    "1111111100001111",
    "1111111011101100",
    "1111111011000001",
    "1111111010010000",
    "1111111001010110",
    "1111111000010110",
    "1111110111010011",
    "1111110110010011",
    "1111110101011101",
    "1111110100111111",
    "1111110101000000",
    "1111110101101010",
    "1111110110111110",
    "1111111001000001",
    "1111111011101001",
    "1111111110101101",
    "1111111110000000",
    "1111111010110110",
    "1111111000000110",
    "1111110101111011",
    "1111110100011110",
    "1111110011101101",
    "1111110011100010",
    "1111110011110101",
    "1111110100011101",
    "1111110101010011",
    "1111110110010100",
    "1111110111011110",
    "1111111000101100",
    "1111111001111101",
    "1111111011010000",
    "1111111100100110",
    "1111111110000001",
    "1111111111100011",
    "1111111110110000",
    "1111111101000111",
    "1111111011100101",
    "1111111010011001",
    "1111111001110000",
    "1111111001101100",
    "1111111010001111",
    "1111111011001100",
    "1111111100011001",
    "1111111101100110",
    "1111111110100111",
    "1111111111011000",
    "1111111111110110",
    "1111111111111001",
    "1111111111111101",
    "1111111111101001",
    "1111111110111101",
    "1111111101110110",
    "1111111100010111",
    "1111111010100100",
    "1111111000101011",
    "1111110110111011",
    "1111110101100100",
    "1111110100110100",
    "1111110100101111",
    "1111110101010111",
    "1111110110100101",
    "1111111000010000",
    "1111111010001110",
    "1111111100010110",
    "1111111110100000",
    "1111111111011010",
    "1111111101100110",
    "1111111100001110",
    "1111111011011100",
    "1111111011010011",
    "1111111011110001",
    "1111111100101101",
    "1111111101110100",
    "1111111110101111",
    "1111111111001000",
    "1111111110110100",
    "1111111101101110",
    "1111111011111100",
    "1111111001101110",
    "1111110111010011",
    "1111110100111100",
    "1111110010110101",
    "1111110001000110",
    "1111101111110110",
    "1111101111001010",
    "1111101111000011",
    "1111101111100010",
    "1111110000100110",
    "1111110010001101",
    "1111110100001100",
    "1111110110010110",
    "1111111000011011",
    "1111111010001101",
    "1111111011100000",
    "1111111100010100",
    "1111111100110010",
    "1111111101001000",
    "1111111101101001",
    "1111111110100001",
    "1111111111110011",
    "1111111110100010",
    "1111111100110000",
    "1111111011000010",
    "1111111001100100",
    "1111111000011001",
    "1111110111100001",
    "1111110110110111",
    "1111110110011001",
    "1111110110001000",
    "1111110110001010",
    "1111110110100111",
    "1111110111100111",
    "1111111001001100",
    "1111111011010010",
    "1111111101101010",
    "1111111111111011",
    "1111111101110101",
    "1111111100010100",
    "1111111011011110",
    "1111111011010110",
    "1111111011110110",
    "1111111100110001",
    "1111111101110100",
    "1111111110110000",
    "1111111111010001",
    "1111111111001100",
    "1111111110010110",
    "1111111100110010",
    "1111111010100100",
    "1111110111111111",
    "1111110101010111",
    "1111110011000001",
    "1111110001010100",
    "1111110000011110",
    "1111110000101000",
    "1111110001101111",
    "1111110011101100",
    "1111110110010000",
    "1111111001001101",
    "1111111100010010",
    "1111111111010001",
    "1111111110000000",
    "1111111011101111",
    "1111111010000100",
    "1111111001000111",
    "1111111001000010",
    "1111111001110110",
    "1111111011100001",
    "1111111101110100",
    "1111111111100110",
    "1111111101010000",
    "1111111011100000",
    "1111111010101001",
    "1111111010101110",
    "1111111011101010",
    "1111111101001001",
    "1111111110110110",
    "1111111111100010",
    "1111111110010100",
    "1111111101100101",
    "1111111101010110",
    "1111111101100011",
    "1111111110001010",
    "1111111111001100",
    "1111111111010001",
    "1111111101010010",
    "1111111010111000",
    "1111111000010000",
    "1111110101101100",
    "1111110011100011",
    "1111110010001001",
    "1111110001101001",
    "1111110010000000",
    "1111110011000011",
    "1111110100011111",
    "1111110101111101",
    "1111110111001000",
    "1111110111111000",
    "1111111000000111",
    "1111110111110111",
    "1111110111010000",
    "1111110110011100",
    "1111110101100000",
    "1111110100100011",
    "1111110011101110",
    "1111110011000011",
    "1111110010101000",
    "1111110010011110",
    "1111110010100011",
    "1111110010110100",
    "1111110011001000",
    "1111110011010111",
    "1111110011011101",
    "1111110011010100",
    "1111110011000000",
    "1111110010100010",
    "1111110010000010",
    "1111110001101000",
    "1111110001011101",
    "1111110001101010",
    "1111110010010110",
    "1111110011100011",
    "1111110101010101",
    "1111110111101010",
    "1111111010011011",
    "1111111101011111",
    "1111111111010100",
    "1111111100010111",
    "1111111001110111",
    "1111111000000101",
    "1111110111001011",
    "1111110111001100",
    "1111111000000100",
    "1111111001101000",
    "1111111011101000",
    "1111111101110001",
    "1111111111110011",
    "1111111110100000",
    "1111111101010010",
    "1111111100100011",
    "1111111100010001",
    "1111111100010011",
    "1111111100100000",
    "1111111100101111",
    "1111111100111001",
    "1111111100110101",
    "1111111100100000",
    "1111111011110110",
    "1111111010110010",
    "1111111001010011",
    "1111110111011010",
    "1111110101001011",
    "1111110010101111",
    "1111110000010010",
    "1111101110000110",
    "1111101100011011",
    "1111101011011111",
    "1111101011011011",
    "1111101100001110",
    "1111101101110110",
    "1111110000001010",
    "1111110010111111",
    "1111110110000111",
    "1111111001010101",
    "1111111100011101",
    "1111111111011000",
    "1111111101111011",
    "1111111011100010",
    "1111111001011011",
    "1111110111101001",
    "1111110110010001",
    "1111110101011000",
    "1111110100111100",
    "1111110100101110",
    "1111110100010101",
    "1111110011000110",
    "1111110000001101",
    "1111101010110011",
    "1111100010000110",
    "1111010101111011",
    "1111000110110010",
    "1110110110011010",
    "1110100111000011",
    "1110011011000100",
    "1110010100000101",
    "1110010010011010",
    "1110010101001000",
    "1110011010010110",
    "1110011111111101",
    "1110100100011010",
    "1110100111000011",
    "1110101000000110",
    "1110101000010101",
    "1110101000100010",
    "1110101001010001",
    "1110101010101011",
    "1110101100100001",
    "1110101110011110",
    "1110110000010101",
    "1110110010010111",
    "1110110101100100",
    "1110111011011110",
    "1111000101100100",
    "1111010100100010",
    "1111101000000110",
    "1111111110111110",
    "1111101000111101",
    "1111010010011010",
    "1110111111100110",
    "1110110001101001",
    "1110101000100010",
    "1110100011010000",
    "1110100000011111",
    "1110011111000111",
    "1110011110010001",
    "1110011101110011",
    "1110011101111011",
    "1110011110111010",
    "1110100000111001",
    "1110100011111110",
    "1110101000101111",
    "1110110000100100",
    "1110111100110010",
    "1111001101110011",
    "1111100010100001",
    "1111111000001010",
    "1111110100110101",
    "1111100111111110",
    "1111100011010011",
    "1111100111000010",
    "1111110001010101",
    "1111111111010110",
    "1111110001110110",
    "1111100100101001",
    "1111011010010110",
    "1111010011011100",
    "1111001111101110",
    "1111001110101011",
    "1111001111100110",
    "1111010001101001",
    "1111010011111110",
    "1111010101110110",
    "1111010110101100",
    "1111010110001011",
    "1111010100100100",
    "1111010010011111",
    "1111010000101001",
    "1111001111100001",
    "1111001111001000",
    "1111001111001101",
    "1111001111011110",
    "1111001111100110",
    "1111001111100100",
    "1111001111010111",
    "1111001111000111",
    "1111001110111000",
    "1111001110110000",
    "1111001110110011",
    "1111001111000000",
    "1111001111100011",
    "1111010000101001",
    "1111010010011100",
    "1111010100111011",
    "1111010111110010",
    "1111011010100010",
    "1111011100100001",
    "1111011101010001",
    "1111011100100011",
    "1111011010100011",
    "1111010111111010",
    "1111010101010111",
    "1111010011100001",
    "1111010010110001",
    "1111010011010111",
    "1111010101010101",
    "1111011000100000",
    "1111011100101010",
    "1111100001010101",
    "1111100110001000",
    "1111101010011111",
    "1111101101110011",
    "1111101111100101",
    "1111101111100110",
    "1111101110000001",
    "1111101011011101",
    "1111101000110100",
    "1111100111001011",
    "1111100111011011",
    "1111101010001001",
    "1111101111011000",
    "1111110110100110",
    "1111111110111110",
    "1111111000011110",
    "1111110000101011",
    "1111101010001000",
    "1111100101000001",
    "1111100001001000",
    "1111011110000010",
    "1111011011001110",
    "1111011000010101",
    "1111010101001101",
    "1111010001111110",
    "1111001110111101",
    "1111001100100101",
    "1111001011001111",
    "1111001011010100",
    "1111001100111000",
    "1111001111111010",
    "1111010100000000",
    "1111011000101111",
    "1111011101100011",
    "1111100001110110",
    "1111100101001011",
    "1111100111001110",
    "1111100111111010",
    "1111100111010100",
    "1111100101101010",
    "1111100011001111",
    "1111100000010010",
    "1111011101001001",
    "1111011001111111",
    "1111010110111111",
    "1111010100010101",
    "1111010010001000",
    "1111010000011100",
    "1111001111010100",
    "1111001110110011",
    "1111001110111010",
    "1111001111100110",
    "1111010000110000",
    "1111010010000110",
    "1111010011011010",
    "1111010100010101",
    "1111010100101110",
    "1111010100011111",
    "1111010011110100",
    "1111010010111110",
    "1111010010010010",
    "1111010010000010",
    "1111010010010000",
    "1111010010111000",
    "1111010011100100",
    "1111010011111100",
    "1111010011101111",
    "1111010010111011",
    "1111010001101100",
    "1111010000011100",
    "1111001111101110",
    "1111001111111101",
    "1111010001010101",
    "1111010011110100",
    "1111010110111111",
    "1111011010010001",
    "1111011100111101",
    "1111011110011111",
    "1111011110101000",
    "1111011101010100",
    "1111011010111010",
    "1111010111110100",
    "1111010100100100",
    "1111010001100001",
    "1111001110110110",
    "1111001100101101",
    "1111001010111100",
    "1111001001100000",
    "1111001000011000",
    "1111000111100111",
    "1111000111010110",
    "1111000111101111",
    "1111001000111010",
    "1111001010111010",
    "1111001101100001",
    "1111010000100011",
    "1111010011100110",
    "1111010110010101",
    "1111011000011010",
    "1111011001100101",
    "1111011001101000",
    "1111011000100000",
    "1111010110001110",
    "1111010010111101",
    "1111001111000101",
    "1111001011001001",
    "1111000111101111",
    "1111000101011111",
    "1111000100110100",
    "1111000101110110",
    "1111001000011011",
    "1111001100000100",
    "1111010000001111",
    "1111010100011000",
    "1111011000001001",
    "1111011011011001",
    "1111011110000101",
    "1111100000010101",
    "1111100010000110",
    "1111100011010111",
    "1111100100000101",
    "1111100100010000",
    "1111100011111011",
    "1111100011001111",
    "1111100010010000",
    "1111100001001000",
    "1111011111111111",
    "1111011110111101",
    "1111011110001100",
    "1111011101111000",
    "1111011110001100",
    "1111011111010111",
    "1111100001100110",
    "1111100100111011",
    "1111101001011000",
    "1111101110111001",
    "1111110101010010",
    "1111111100010111",
    "1111111100001110",
    "1111110100110111",
    "1111101101111010",
    "1111100111100111",
    "1111100010001101",
    "1111011101111000",
    "1111011010110010",
    "1111011001000111",
    "1111011000111110",
    "1111011010011001",
    "1111011101010110",
    "1111100001100110",
    "1111100110110110",
    "1111101100101100",
    "1111110010101010",
    "1111111000001101",
    "1111111100110111",
    "1111111111101001",
    "1111111101100010",
    "1111111100100111",
    "1111111100100011",
    "1111111101000110",
    "1111111110000010",
    "1111111111010101",
    "1111111110111111",
    "1111111101001001",
    "1111111011100000",
    "1111111010011110",
    "1111111010010011",
    "1111111010111111",
    "1111111100010100",
    "1111111110000101",
    "1111111111110110",
    "1111111101101011",
    "1111111011011111",
    "1111111001101001",
    "1111111000100101",
    "1111111000101111",
    "1111111010010111",
    "1111111101010111",
    "1111111110101000",
    "1111111010001000",
    "1111110101100100",
    "1111110001000110",
    "1111101100110011",
    "1111101000101001",
    "1111100100101001",
    "1111100000111001",
    "1111011101100011",
    "1111011010110111",
    "1111011001000110",
    "1111011000011011",
    "1111011000101010",
    "1111011001010011",
    "1111011001011101",
    "1111011000010101",
    "1111010101011011",
    "1111010001000000",
    "1111001100000010",
    "1111000111110111",
    "1111000101101001",
    "1111000101110111",
    "1111001000000110",
    "1111001011010001",
    "1111001110000101",
    "1111001111101001",
    "1111001111101000",
    "1111001110011001",
    "1111001100101011",
    "1111001011010001",
    "1111001010110010",
    "1111001011011110",
    "1111001101010100",
    "1111010000000010",
    "1111010011010000",
    "1111010110101101",
    "1111011001111101",
    "1111011100101110",
    "1111011110101001",
    "1111011111011100",
    "1111011110110101",
    "1111011100101101",
    "1111011001000001",
    "1111010100000101",
    "1111001110010111",
    "1111001000101100",
    "1111000011111001",
    "1111000000111000",
    "1111000000011110",
    "1111000011001111",
    "1111001001010110",
    "1111010010011111",
    "1111011101101011",
    "1111101001011011",
    "1111110011111101",
    "1111111011100100",
    "1111111110101111",
    "1111111100010101",
    "1111110011001110",
    "1111100010101111",
    "1111001011011001",
    "1110101111010010",
    "1110010010000000",
    "1101110111110010",
    "1101100100011101",
    "1101011010011000",
    "1101011001101101",
    "1101100000001010",
    "1101101010010001",
    "1101110100011111",
    "1101111100010110",
    "1110000000111110",
    "1110000010110100",
    "1110000011001011",
    "1110000011010011",
    "1110000100000000",
    "1110000101010000",
    "1110000110100010",
    "1110000111001101",
    "1110000110110010",
    "1110000101010111",
    "1110000011000110",
    "1110000000011100",
    "1101111101101000",
    "1101111011000111",
    "1101111001100010",
    "1101111010110000",
    "1110000010000000",
    "1110010010000010",
    "1110101011101101",
    "1111001101000010",
    "1111110001001100",
    "1111101101101101",
    "1111010101000001",
    "1111000111100010",
    "1111000100001101",
    "1111000111010011",
    "1111001100010100",
    "1111001111101110",
    "1111010000000111",
    "1111001101111011",
    "1111001010100101",
    "1111000111011011",
    "1111000100111100",
    "1111000010100111",
    "1110111111100110",
    "1110111011001111",
    "1110110101100101",
    "1110101111010010",
    "1110101001011001",
    "1110100100101001",
    "1110100001000101",
    "1110011110011001",
    "1110011100001010",
    "1110011010010001",
    "1110011000110101",
    "1110011000000001",
    "1110010111111111",
    "1110011000110111",
    "1110011010100011",
    "1110011101001010",
    "1110100000101110",
    "1110100101011000",
    "1110101011001001",
    "1110110001110100",
    "1110111010001111",
    "1111000110100111",
    "1111011000111111",
    "1111110001111100",
    "1111110000101111",
    "1111010011101110",
    "1110111100001001",
    "1110101110001111",
    "1110101011110000",
    "1110110010111000",
    "1110111111010111",
    "1111001100100001",
    "1111010111000011",
    "1111011110010010",
    "1111100011110011",
    "1111101001111111",
    "1111110011001101",
    "1111111111101011",
    "1111101111110100",
    "1111011111011100",
    "1111010001001000",
    "1111000110111001",
    "1111000001010101",
    "1110111111110000",
    "1111000000110011",
    "1111000011000110",
    "1111000101110100",
    "1111001000010101",
    "1111001010001100",
    "1111001011011001",
    "1111001100001110",
    "1111001101001010",
    "1111001110110011",
    "1111010001010101",
    "1111010100110110",
    "1111011000111111",
    "1111011101011011",
    "1111100001101011",
    "1111100101011111",
    "1111101000111100",
    "1111101100011010",
    "1111110000011001",
    "1111110101001111",
    "1111111010111110",
    "1111111110110000",
    "1111111000100110",
    "1111110011001000",
    "1111101110011101",
    "1111101010010100",
    "1111100110001000",
    "1111100001100001",
    "1111011100100001",
    "1111010111101010",
    "1111010011100001",
    "1111010000011100",
    "1111001110011100",
    "1111001101001110",
    "1111001100011001",
    "1111001011101101",
    "1111001011001010",
    "1111001011001001",
    "1111001100001100",
    "1111001110101101",
    "1111010010100001",
    "1111010111000011",
    "1111011011011001",
    "1111011110110011",
    "1111100000110101",
    "1111100001011111",
    "1111100001011001",
    "1111100001011100",
    "1111100010010101",
    "1111100100010011",
    "1111100111000111",
    "1111101010000000",
    "1111101100001010",
    "1111101100111101",
    "1111101100001001",
    "1111101001111011",
    "1111100110111010",
    "1111100011110100",
    "1111100001010010",
    "1111011111101001",
    "1111011111000100",
    "1111011111100011",
    "1111100001001101",
    "1111100100001101",
    "1111101000110001",
    "1111101111000011",
    "1111110110111110",
    "1111111111101111",
    "1111110101110100",
    "1111101100000001",
    "1111100011001111",
    "1111011100001110",
    "1111010111100010",
    "1111010101011000",
    "1111010101101110",
    "1111011000001000",
    "1111011100000101",
    "1111100000111110",
    "1111100110001000",
    "1111101010111001",
    "1111101110111000",
    "1111110001110010",
    "1111110011100001",
    "1111110100001110",
    "1111110100001010",
    "1111110011101111",
    "1111110011011010",
    "1111110011100001",
    "1111110100001010",
    "1111110101001010",
    "1111110110001110",
    "1111110111000010",
    "1111110111011001",
    "1111110111011011",
    "1111110111011011",
    "1111110111110100",
    "1111111000110001",
    "1111111010010001",
    "1111111011111110",
    "1111111101010111",
    "1111111101111101",
    "1111111101011111",
    "1111111100000001",
    "1111111001111000",
    "1111110111100101",
    "1111110101101110",
    "1111110100101000",
    "1111110100011010",
    "1111110100110100",
    "1111110101010110",
    "1111110101010101",
    "1111110100010011",
    "1111110010001001",
    "1111101111001011",
    "1111101100000001",
    "1111101001011001",
    "1111100111111110",
    "1111101000000001",
    "1111101001100110",
    "1111101100010111",
    "1111101111101011",
    "1111110010101101",
    "1111110100101001",
    "1111110100110101",
    "1111110011000010",
    "1111101111100010",
    "1111101011000100",
    "1111100110100101",
    "1111100010111000",
    "1111100000010111",
    "1111011111000100",
    "1111011110101000",
    "1111011110101000",
    "1111011110101000",
    "1111011110010010",
    "1111011101011110",
    "1111011100001001",
    "1111011010011110",
    "1111011000110010",
    "1111010111011010",
    "1111010110100101",
    "1111010110010010",
    "1111010110001001",
    "1111010101101110",
    "1111010100011101",
    "1111010001111110",
    "1111001110010010",
    "1111001001100101",
    "1111000100010101",
    "1110111111000100",
    "1110111010010110",
    "1110110110100101",
    "1110110100000011",
    "1110110010101011",
    "1110110010001011",
    "1110110010001101",
    "1110110010100010",
    "1110110011010000",
    "1110110100101100",
    "1110110111010101",
    "1110111011011001",
    "1111000000110101",
    "1111000111000100",
    "1111001101100011",
    "1111010011101010",
    "1111011001001110",
    "1111011110010001",
    "1111100010111000",
    "1111100111000001",
    "1111101010011010",
    "1111101100101101",
    "1111101101101001",
    "1111101101001111",
    "1111101011110110",
    "1111101001111111",
    "1111101000000101",
    "1111100110001011",
    "1111100100000101",
    "1111100001011010",
    "1111011101111111",
    "1111011010001001",
    "1111010110101100",
    "1111010100110100",
    "1111010101101100",
    "1111011001110111",
    "1111100001000010",
    "1111101001111111",
    "1111110011000000",
    "1111111010010111",
    "1111111110111011",
    "1111111111011011",
    "1111111111111001",
    "1111111110001011",
    "1111111100011101",
    "1111111011010011",
    "1111111010011111",
    "1111111001010011",
    "1111110110111000",
    "1111110010110010",
    "1111101101001110",
    "1111100111000010",
    "1111100001011001",
    "1111011101010110",
    "1111011011100000",
    "1111011011111010",
    "1111011110000101",
    "1111100001010000",
    "1111100100101110",
    "1111100111101100",
    "1111101001101011",
    "1111101010010001",
    "1111101001010011",
    "1111100110110011",
    "1111100011001011",
    "1111011111000000",
    "1111011011000111",
    "1111011000001000",
    "1111010110010101",
    "1111010101011111",
    "1111010100111001",
    "1111010011101010",
    "1111010001010000",
    "1111001101101011",
    "1111001001101000",
    "1111000110010101",
    "1111000101000001",
    "1111000110011111",
    "1111001010110100",
    "1111010001010101",
    "1111011001000110",
    "1111100000111101",
    "1111101000010101",
    "1111101111000110",
    "1111110101100100",
    "1111111100001001",
    "1111111100111010",
    "1111110101111000",
    "1111101111011000",
    "1111101010010110",
    "1111100111101011",
    "1111100111111010",
    "1111101011000000",
    "1111110000010000",
    "1111110110010111",
    "1111111011110111",
    "1111111111010010",
    "1111111111101001",
    "1111111100100110",
    "1111110110100001",
    "1111101110011110",
    "1111100101111100",
    "1111011110100110",
    "1111011001111100",
    "1111011001000100",
    "1111011100011001",
    "1111100011100111",
    "1111101101100011",
    "1111111000100011",
    "1111111101010001",
    "1111110101110001",
    "1111110010010000",
    "1111110011011111",
    "1111111001101110",
    "1111111011011011",
    "1111101101000001",
    "1111011100110000",
    "1111001100110010",
    "1110111111010111",
    "1110110110100010",
    "1110110011101110",
    "1110110111101101",
    "1111000010100010",
    "1111010011011010",
    "1111101000101000",
    "1111111111100111",
    "1111101010100100",
    "1111011000110100",
    "1111001101000000",
    "1111000111110111",
    "1111001000110111",
    "1111001110110000",
    "1111011000001100",
    "1111100100001110",
    "1111110010100011",
    "1111111100111100",
    "1111101010110001",
    "1111011000000001",
    "1111000110010101",
    "1110110111100010",
    "1110101100110101",
    "1110100110011010",
    "1110100011001101",
    "1110100001011111",
    "1110011111101011",
    "1110011101001110",
    "1110011010100101",
    "1110011000110111",
    "1110011000111111",
    "1110011011000100",
    "1110011110001111",
    "1110100001000000",
    "1110100001111001",
    "1110100000000101",
    "1110011011100110",
    "1110010101001101",
    "1110001110001001",
    "1110000111100000",
    "1110000010001011",
    "1101111110100110",
    "1101111100110111",
    "1101111100111000",
    "1101111110100011",
    "1110000001100111",
    "1110000101110001",
    "1110001010100101",
    "1110001111100100",
    "1110010100011010",
    "1110011001100111",
    "1110100001000011",
    "1110101101011100",
    "1111000000111101",
    "1111011011101101",
    "1111111011001010",
    "1111100101011010",
    "1111001011011110",
    "1110111011001111",
    "1110110110001011",
    "1110111010011001",
    "1111000011111001",
    "1111001110000000",
    "1111010101001001",
    "1111010111110100",
    "1111010110001110",
    "1111010001110001",
    "1111001100000010",
    "1111000110001000",
    "1111000000011100",
    "1110111011000010",
    "1110110101111001",
    "1110110001010000",
    "1110101101110010",
    "1110101011111100",
    "1110101011110111",
    "1110101101001110",
    "1110101111010001",
    "1110110001010111",
    "1110110011001010",
    "1110110100011100",
    "1110110101001101",
    "1110110101100010",
    "1110110101011111",
    "1110110101010000",
    "1110110101110110",
    "1110111001111111",
    "1111000101001001",
    "1111011001100000",
    "1111110110011101",
    "1111100111111001",
    "1111000111110010",
    "1110101111011001",
    "1110100011001111",
    "1110100011111100",
    "1110101110010010",
    "1110111100111100",
    "1111001010110000",
    "1111010100101010",
    "1111011010011101",
    "1111011101101101",
    "1111100000110110",
    "1111100101111100",
    "1111101101100100",
    "1111110111001000",
    "1111111110100000",
    "1111110100110100",
    "1111101100101011",
    "1111100110011011",
    "1111100010001010",
    "1111100000000010",
    "1111100000010101",
    "1111100011000110",
    "1111100111101010",
    "1111101100110101",
    "1111110001011110",
    "1111110100100101",
    "1111110101111000",
    "1111110101101010",
    "1111110100101001",
    "1111110011110000",
    "1111110011110100",
    "1111110101010011",
    "1111111000010110",
    "1111111100111010",
    "1111111101010001",
    "1111110110101111",
    "1111110000000101",
    "1111101001111111",
    "1111100101000001",
    "1111100001100110",
    "1111011111110011",
    "1111011111010110",
    "1111011111100110",
    "1111011111110110",
    "1111011111011100",
    "1111011110000000",
    "1111011011011011",
    "1111010111110010",
    "1111010011010111",
    "1111001110011110",
    "1111001001011110",
    "1111000100110001",
    "1111000000100011",
    "1110111100111111",
    "1110111010010011",
    "1110111000110111",
    "1110111001000001",
    "1110111010110101",
    "1110111101111011",
    "1111000001100110",
    "1111000101000011",
    "1111000111101000",
    "1111001001001100",
    "1111001001111001",
    "1111001010001110",
    "1111001010101000",
    "1111001011011000",
    "1111001100100000",
    "1111001101111111",
    "1111001111110000",
    "1111010001101011",
    "1111010011011010",
    "1111010100101001",
    "1111010100110111",
    "1111010011111001",
    "1111010001101100",
    "1111001110101101",
    "1111001011100101",
    "1111001001001100",
    "1111001000011010",
    "1111001001101101",
    "1111001101010010",
    "1111010010111001",
    "1111011001110101",
    "1111100001001010",
    "1111100111110111",
    "1111101101001110",
    "1111110000110011",
    "1111110010101100",
    "1111110011010101",
    "1111110011010101",
    "1111110011010101",
    "1111110011110000",
    "1111110100110001",
    "1111110110001111",
    "1111110111110100",
    "1111111001000010",
    "1111111001100010",
    "1111111001000110",
    "1111110111110111",
    "1111110110010010",
    "1111110101000000",
    "1111110100110000",
    "1111110101110101",
    "1111111000000100",
    "1111111010110000",
    "1111111100111100",
    "1111111101101101",
    "1111111100100010",
    "1111111001100010",
    "1111110101011001",
    "1111110001000001",
    "1111101101001101",
    "1111101010011001",
    "1111101000100001",
    "1111100111001101",
    "1111100110000011",
    "1111100100110110",
    "1111100011101100",
    "1111100010111101",
    "1111100011000001",
    "1111100100010010",
    "1111100110110011",
    "1111101010011010",
    "1111101110101111",
    "1111110011010000",
    "1111110111100010",
    "1111111011010010",
    "1111111110010000",
    "1111111111100011",
    "1111111110010101",
    "1111111110000101",
    "1111111110101111",
    "1111111111110110",
    "1111111110010001",
    "1111111101000110",
    "1111111100111101",
    "1111111110010100",
    "1111111110101101",
    "1111111010100100",
    "1111110101111001",
    "1111110001011101",
    "1111101101110011",
    "1111101011000111",
    "1111101001010000",
    "1111100111110101",
    "1111100110011110",
    "1111100101000000",
    "1111100011100110",
    "1111100010100111",
    "1111100010011101",
    "1111100011010011",
    "1111100100111011",
    "1111100110110101",
    "1111101000010100",
    "1111101000111000",
    "1111101000010101",
    "1111100110111101",
    "1111100101010101",
    "1111100100000101",
    "1111100011100111",
    "1111100011111110",
    "1111100100110001",
    "1111100101010101",
    "1111100100111110",
    "1111100011010101",
    "1111100000010101",
    "1111011100001110",
    "1111010111011011",
    "1111010010011101",
    "1111001101101101",
    "1111001001011101",
    "1111000110000001",
    "1111000011101110",
    "1111000010110001",
    "1111000011010011",
    "1111000101001110",
    "1111001000001000",
    "1111001011011110",
    "1111001110101110",
    "1111010001100100",
    "1111010011111100",
    "1111010110001011",
    "1111011000100101",
    "1111011011010110",
    "1111011110010001",
    "1111100000111001",
    "1111100010100010",
    "1111100010101001",
    "1111100001000000",
    "1111011101110011",
    "1111011001110100",
    "1111010101110111",
    "1111010010111001",
    "1111010001011111",
    "1111010001101110",
    "1111010011011010",
    "1111010101111100",
    "1111011000110100",
    "1111011011100001",
    "1111011101111101",
    "1111100000001101",
    "1111100010100001",
    "1111100101000011",
    "1111100111111000",
    "1111101010110011",
    "1111101101011110",
    "1111101111011111",
    "1111110000011110",
    "1111110000010001",
    "1111101110111100",
    "1111101100110110",
    "1111101010100011",
    "1111101000101100",
    "1111100111101101",
    "1111100111110000",
    "1111101000100011",
    "1111101001011110",
    "1111101001110100",
    "1111101000111110",
    "1111100110101001",
    "1111100011000101",
    "1111011110110000",
    "1111011010100000",
    "1111010111001000",
    "1111010101001011",
    "1111010100111110",
    "1111010110011010",
    "1111011000111111",
    "1111011011111101",
    "1111011110011100",
    "1111011111011111",
    "1111011110011111",
    "1111011011000110",
    "1111010101011000",
    "1111001101111011",
    "1111000101100111",
    "1110111101100100",
    "1110110111000011",
    "1110110011000101",
    "1110110010011100",
    "1110110101011000",
    "1110111011100110",
    "1111000100010000",
    "1111001110000111",
    "1111010111110100",
    "1111100000000101",
    "1111100101111110",
    "1111101001000010",
    "1111101001001100",
    "1111100110110101",
    "1111100010100100",
    "1111011101010100",
    "1111011000001011",
    "1111010100010101",
    "1111010010111110",
    "1111010101000110",
    "1111011011001100",
    "1111100100111110",
    "1111110001010100",
    "1111111110010111",
    "1111110110000000",
    "1111101101110101",
    "1111101010011100",
    "1111101100011100",
    "1111110011101001",
    "1111111111010000",
    "1111110010000110",
    "1111100010011001",
    "1111010011101010",
    "1111000111111110",
    "1111000001000000",
    "1110111111111101",
    "1111000101010111",
    "1111010000111101",
    "1111100001101001",
    "1111110101011101",
    "1111110110000111",
    "1111100011110100",
    "1111010101110110",
    "1111001101100000",
    "1111001010111101",
    "1111001101101000",
    "1111010100011111",
    "1111011110101110",
    "1111101011101000",
    "1111111010100100",
    "1111110101011101",
    "1111100110000001",
    "1111011000110101",
    "1111001111011111",
    "1111001011000001",
    "1111001011011101",
    "1111001111101110",
    "1111010110000001",
    "1111011100001100",
    "1111100000100001",
    "1111100010001011",
    "1111100001010010",
    "1111011110110101",
    "1111011100000111",
    "1111011010100010",
    "1111011011010100",
    "1111011111011110",
    "1111100111111010",
    "1111110101000100",
    "1111111001101010",
    "1111100110001011",
    "1111010011000101",
    "1111000011001000",
    "1110111000010001",
    "1110110011001111",
    "1110110011000110",
    "1110110101111001",
    "1110111001001011",
    "1110111011000001",
    "1110111010011011",
    "1110110111100011",
    "1110110011001010",
    "1110101110010100",
    "1110101001110111",
    "1110100110010011",
    "1110100011100100",
    "1110100001100010",
    "1110100000000010",
    "1110011111000000",
    "1110011110010111",
    "1110011110000111",
    "1110011110000010",
    "1110011101111101",
    "1110011101111010",
    "1110011110000101",
    "1110011110101110",
    "1110100000100111",
    "1110100101101010",
    "1110110000010111",
    "1111000010011100",
    "1111011011101000",
    "1111111001001011",
    "1111101001011111",
    "1111010001010100",
    "1111000001111110",
    "1110111100011011",
    "1110111110101001",
    "1111000100111110",
    "1111001011011001",
    "1111001111000111",
    "1111001111010100",
    "1111001100100011",
    "1111001000010001",
    "1111000100000001",
    "1111000000110011",
    "1110111110110110",
    "1110111110000010",
    "1110111101110111",
    "1110111110000010",
    "1110111110100001",
    "1110111111001101",
    "1110111111110001",
    "1110111111011111",
    "1110111101110000",
    "1110111010011000",
    "1110110101101110",
    "1110110000100001",
    "1110101011101111",
    "1110101000010110",
    "1110100111001110",
    "1110101000111010",
    "1110101101100100",
    "1110110100111001",
    "1110111110011100",
    "1111001010011011",
    "1111011001111100",
    "1111101101101110",
    "1111111010100110",
    "1111100001001010",
    "1111001001011101",
    "1110110111000110",
    "1110101100110010",
    "1110101011000010",
    "1110101111110011",
    "1110110111100000",
    "1110111110101101",
    "1111000011000110",
    "1111000100011000",
    "1111000011110100",
    "1111000011011010",
    "1111000101010010",
    "1111001010100110",
    "1111010011001101",
    "1111011101110111",
    "1111101000110110",
    "1111110010101011",
    "1111111010100001",
    "1111111111110101",
    "1111111100011001",
    "1111111010111101",
    "1111111011001101",
    "1111111100110010",
    "1111111111000101",
    "1111111110010110",
    "1111111100000011",
    "1111111010001100",
    "1111111000110010",
    "1111110111101101",
    "1111110110101111",
    "1111110101101110",
    "1111110100101001",
    "1111110011100011",
    "1111110010100000",
    "1111110001011000",
    "1111101111111010",
    "1111101101101000",
    "1111101010000110",
    "1111100101001001",
    "1111011111000101",
    "1111011000101100",
    "1111010010110100",
    "1111001110000100",
    "1111001010011001",
    "1111000111011000",
    "1111000100001000",
    "1110111111111101",
    "1110111010100010",
    "1110110100000101",
    "1110101101010110",
    "1110100111010110",
    "1110100011000110",
    "1110100001010100",
    "1110100010000101",
    "1110100100111110",
    "1110101001001100",
    "1110101101110111",
    "1110110010001101",
    "1110110101101010",
    "1110111000001001",
    "1110111001101101",
    "1110111010101011",
    "1110111011001111",
    "1110111011100001",
    "1110111011100011",
    "1110111011100000",
    "1110111011100110",
    "1110111100010110",
    "1110111110001001",
    "1111000001001100",
    "1111000101010010",
    "1111001001110100",
    "1111001101111000",
    "1111010000101110",
    "1111010001111101",
    "1111010001101001",
    "1111010000010111",
    "1111001110110101",
    "1111001101101110",
    "1111001101011110",
    "1111001110001100",
    "1111001111101100",
    "1111010001111000",
    "1111010100101001",
    "1111010111111111",
    "1111011100000101",
    "1111100000110011",
    "1111100101110110",
    "1111101010100001",
    "1111101110001100",
    "1111110000011011",
    "1111110001010001",
    "1111110001001110",
    "1111110001001010",
    "1111110001111000",
    "1111110011110010",
    "1111110110110101",
    "1111111010011101",
    "1111111101111001",
    "1111111111100001",
    "1111111110010000",
    "1111111110010101",
    "1111111111100010",
    "1111111110011110",
    "1111111100001010",
    "1111111001110011",
    "1111110111101000",
    "1111110101101110",
    "1111110100001010",
    "1111110010110101",
    "1111110001101010",
    "1111110000100010",
    "1111101111010001",
    "1111101101110111",
    "1111101100011011",
    "1111101011001100",
    "1111101010100010",
    "1111101010110000",
    "1111101100000110",
    "1111101110100101",
    "1111110001111010",
    "1111110101100100",
    "1111111000111011",
    "1111111011011101",
    "1111111100110111",
    "1111111101010010",
    "1111111101001010",
    "1111111101000111",
    "1111111101110100",
    "1111111111101000",
    "1111111101011001",
    "1111111001101100",
    "1111110101110110",
    "1111110010011111",
    "1111110000001010",
    "1111101111000101",
    "1111101110111110",
    "1111101111010110",
    "1111101111011101",
    "1111101110110010",
    "1111101101001001",
    "1111101010110101",
    "1111101000011111",
    "1111100110111100",
    "1111100110101111",
    "1111100111111101",
    "1111101010001001",
    "1111101100011111",
    "1111101110001001",
    "1111101110100001",
    "1111101101011110",
    "1111101011010011",
    "1111101000100111",
    "1111100110001011",
    "1111100100101001",
    "1111100100011000",
    "1111100101010101",
    "1111100111000101",
    "1111101001000000",
    "1111101010010111",
    "1111101010100010",
    "1111101001001111",
    "1111100110100011",
    "1111100010111000",
    "1111011110110101",
    "1111011010111100",
    "1111010111101100",
    "1111010101010010",
    "1111010011101110",
    "1111010010110110",
    "1111010010011101",
    "1111010010011010",
    "1111010010100110",
    "1111010010111110",
    "1111010011100001",
    "1111010100010000",
    "1111010101011000",
    "1111010111000011",
    "1111011001100000",
    "1111011100110111",
    "1111100001001010",
    "1111100110010000",
    "1111101011110110",
    "1111110001100101",
    "1111110111000100",
    "1111111011111101",
    "1111111111111011",
    "1111111100101111",
    "1111111010011011",
    "1111111000111011",
    "1111111000001111",
    "1111111000011000",
    "1111111001100101",
    "1111111100000111",
    "1111111111101010",
    "1111111001101101",
    "1111110001111111",
    "1111101000100111",
    "1111011101110111",
    "1111010010001010",
    "1111000110001110",
    "1110111010111100",
    "1110110001010100",
    "1110101010001001",
    "1110100101101111",
    "1110100011111011",
    "1110100100000000",
    "1110100100110111",
    "1110100101011101",
    "1110100100111011",
    "1110100010111001",
    "1110011111011100",
    "1110011011000111",
    "1110010110100111",
    "1110010010110011",
    "1110010000010111",
    "1110001111110110",
    "1110010001101001",
    "1110010101111011",
    "1110011100110011",
    "1110100110010011",
    "1110110001111001",
    "1110111110101110",
    "1111001011010011",
    "1111010110000100",
    "1111011101101110",
    "1111100001100010",
    "1111100001101100",
    "1111011111010110",
    "1111011100001100",
    "1111011010001100",
    "1111011010111100",
    "1111011111001100",
    "1111100110110010",
    "1111110000100110",
    "1111111011000000",
    "1111111011110110",
    "1111110101100001",
    "1111110010111011",
    "1111110100011000",
    "1111111001110010",
    "1111111101001000",
    "1111110000110011",
    "1111100001111101",
    "1111010001111101",
    "1111000010101100",
    "1110110110010110",
    "1110101110110101",
    "1110101101011011",
    "1110110010011001",
    "1110111101001110",
    "1111001100110101",
    "1111011111110110",
    "1111110100100111",
    "1111110110110101",
    "1111100100110011",
    "1111010111011010",
    "1111010000011010",
    "1111010000110000",
    "1111011000010101",
    "1111100101111100",
    "1111110111100001",
    "1111110101101000",
    "1111100100010011",
    "1111010110110010",
    "1111001110100100",
    "1111001100010111",
    "1111010000000000",
    "1111011000110010",
    "1111100101100111",
    "1111110101000110",
    "1111111010010010",
    "1111101010010010",
    "1111011100100000",
    "1111010010001010",
    "1111001011111100",
    "1111001001111001",
    "1111001011100000",
    "1111001111110001",
    "1111010101100100",
    "1111011011101010",
    "1111100000111101",
    "1111100100101110",
    "1111100110100111",
    "1111100110101101",
    "1111100101100000",
    "1111100011111000",
    "1111100010111101",
    "1111100100000001",
    "1111101000000010",
    "1111101111001110",
    "1111111000111001",
    "1111111100011011",
    "1111110010101011",
    "1111101011010110",
    "1111100111001110",
    "1111100110001000",
    "1111100111010110",
    "1111101001111011",
    "1111101101011000",
    "1111110001111001",
    "1111111000001101",
    "1111111110101110",
    "1111110010011110",
    "1111100011010111",
    "1111010010110110",
    "1111000011001000",
    "1110110110011010",
    "1110101110000010",
    "1110101010000111",
    "1110101001100000",
    "1110101010100000",
    "1110101011100000",
    "1110101011101000",
    "1110101010110010",
    "1110101001100000",
    "1110101000011101",
    "1110101000000100",
    "1110101000010001",
    "1110101000110010",
    "1110101001001001",
    "1110101001000111",
    "1110101000110000",
    "1110101000010011",
    "1110100111111001",
    "1110100111101000",
    "1110100111010011",
    "1110100110100101",
    "1110100101010011",
    "1110100011011010",
    "1110100001001101",
    "1110011111001000",
    "1110011101101000",
    "1110011101000101",
    "1110011101111000",
    "1110100000001111",
    "1110100100011100",
    "1110101010101010",
    "1110110010111110",
    "1110111101010010",
    "1111001001010001",
    "1111010110011111",
    "1111100100011000",
    "1111110010101101",
    "1111111110011100",
    "1111101111001000",
    "1111011111101000",
    "1111010000110011",
    "1111000011111011",
    "1110111010011001",
    "1110110101000000",
    "1110110011100110",
    "1110110101000000",
    "1110110111011000",
    "1110111000111110",
    "1110111000100101",
    "1110110110000000",
    "1110110001111011",
    "1110101101100000",
    "1110101001111001",
    "1110100111110111",
    "1110100111100011",
    "1110101000101000",
    "1110101010100000",
    "1110101100100110",
    "1110101110011110",
    "1110101111110110",
    "1110110000100011",
    "1110110000011001",
    "1110101111010110",
    "1110101101100100",
    "1110101011110111",
    "1110101100010001",
    "1110110010000010",
    "1110111111101100",
    "1111010101101110",
    "1111110001101010",
    "1111110001001011",
    "1111011000010110",
    "1111001000011000",
    "1111000011010111",
    "1111000111111100",
    "1111010010100001",
    "1111011111000010",
    "1111101010011111",
    "1111110011110000",
    "1111111011010010",
    "1111111101110010",
    "1111110110100000",
    "1111101110100111",
    "1111100110110000",
    "1111011111111000",
    "1111011010110101",
    "1111010111111111",
    "1111010111000100",
    "1111010111100011",
    "1111011001000100",
    "1111011011100101",
    "1111011111001010",
    "1111100011100010",
    "1111101000001001",
    "1111101100001110",
    "1111101111000111",
    "1111110000011001",
    "1111110000000100",
    "1111101110011011",
    "1111101100000000",
    "1111101001010011",
    "1111100110101110",
    "1111100100011111",
    "1111100010110110",
    "1111100010000110",
    "1111100010110001",
    "1111100101011000",
    "1111101010011000",
    "1111110001111010",
    "1111111011100000",
    "1111111001110000",
    "1111101111001100",
    "1111100101111001",
    "1111011110100110",
    "1111011001100111",
    "1111010110111100",
    "1111010110010010",
    "1111010111000100",
    "1111011000011110",
    "1111011001011011",
    "1111011000101111",
    "1111010101100010",
    "1111001111011010",
    "1111000110100101",
    "1110111011110101",
    "1110110000010100",
    "1110100101010010",
    "1110011011100110",
    "1110010011100111",
    "1110001101000111",
    "1110000111101010",
    "1110000010110100",
    "1101111110011100",
    "1101111010101011",
    "1101111000001100",
    "1101110111101101",
    "1101111001110111",
    "1101111111000000",
    "1110000111001001",
    "1110010001110100",
    "1110011110011011",
    "1110101100000010",
    "1110111001110101",
    "1111000111001001",
    "1111010011100010",
    "1111011111000000",
    "1111101001101110",
    "1111110100000001",
    "1111111110000011",
    "1111111000001000",
    "1111101110110000",
    "1111100101111110",
    "1111011101111011",
    "1111010110100101",
    "1111001111101100",
    "1111001001001001",
    "1111000010110110",
    "1110111100111000",
    "1110110111100101",
    "1110110011010000",
    "1110110000001101",
    "1110101110101000",
    "1110101110100011",
    "1110101111111101",
    "1110110010110100",
    "1110110111001001",
    "1110111100111111",
    "1111000100010011",
    "1111001100111111",
    "1111010110111011",
    "1111100001111000",
    "1111101101101100",
    "1111111010000110",
    "1111111001001100",
    "1111101100101110",
    "1111100001001000",
    "1111010111000110",
    "1111001111001100",
    "1111001001110101",
    "1111000111000110",
    "1111000110101101",
    "1111001000010011",
    "1111001011010011",
    "1111001111001100",
    "1111010011100010",
    "1111011000000011",
    "1111011100011011",
    "1111100000100100",
    "1111100100011101",
    "1111101000010001",
    "1111101100000101",
    "1111110000000100",
    "1111110100001110",
    "1111111000011010",
    "1111111100010100",
    "1111111111100101",
    "1111111110001000",
    "1111111101001101",
    "1111111101110001",
    "1111111111101110",
    "1111111101010110",
    "1111111010000111",
    "1111110111010101",
    "1111110101100111",
    "1111110101010010",
    "1111110110001101",
    "1111110111110001",
    "1111111001001010",
    "1111111001110010",
    "1111111001011001",
    "1111111000001110",
    "1111110110110100",
    "1111110101110111",
    "1111110101111001",
    "1111110111001011",
    "1111111001011101",
    "1111111100001111",
    "1111111110110101",
    "1111111111010110",
    "1111111110101110",
    "1111111111010001",
    "1111111111010101",
    "1111111101101010",
    "1111111100001101",
    "1111111011010011",
    "1111111011001001",
    "1111111011110001",
    "1111111101001001",
    "1111111111001000",
    "1111111110011111",
    "1111111100001001",
    "1111111010010000",
    "1111111001001010",
    "1111111001000000",
    "1111111001101100",
    "1111111010111101",
    "1111111100010101",
    "1111111101011010",
    "1111111101111010",
    "1111111101101010",
    "1111111100101010",
    "1111111011000000",
    "1111111000101111",
    "1111110110000011",
    "1111110011001101",
    "1111110000100101",
    "1111101110101000",
    "1111101101110101",
    "1111101110100100",
    "1111110001000100",
    "1111110101010001",
    "1111111010101010",
    "1111111111100010",
    "1111111010011011",
    "1111110111000010",
    "1111110110001100",
    "1111111000011100",
    "1111111101101111",
    "1111111010100111",
    "1111110001110110",
    "1111101001011111",
    "1111100011000011",
    "1111011111101100",
    "1111100000000011",
    "1111100100000000",
    "1111101010101000",
    "1111110010100011",
    "1111111010010000",
    "1111111111100100",
    "1111111011111001",
    "1111111010111110",
    "1111111100101001",
    "1111111111100100",
    "1111111010011100",
    "1111110100101011",
    "1111101111000101",
    "1111101010011101",
    "1111100111101100",
    "1111100111100001",
    "1111101010010010",
    "1111101111110101",
    "1111110111010101",
    "1111111111011110",
    "1111111001001100",
    "1111110100000010",
    "1111110001111100",
    "1111110011010111",
    "1111111000010010",
    "1111111111100010",
    "1111110100110000",
    "1111101000010010",
    "1111011011100001",
    "1111010000010001",
    "1111001000010110",
    "1111000101010010",
    "1111000111110101",
    "1111001111101100",
    "1111011011011101",
    "1111101000111100",
    "1111110101101110",
    "1111111111101001",
    "1111111010100101",
    "1111111001100000",
    "1111111100110011",
    "1111111100000010",
    "1111110001101011",
    "1111100100110111",
    "1111010110110001",
    "1111001000111110",
    "1110111101010001",
    "1110110101011011",
    "1110110010101100",
    "1110110101100101",
    "1110111101101110",
    "1111001010000100",
    "1111011001001001",
    "1111101001001010",
    "1111111000001100",
    "1111111011100010",
    "1111110011101010",
    "1111110001001010",
    "1111110100001001",
    "1111111011111100",
    "1111111000110011",
    "1111101011111010",
    "1111011111000010",
    "1111010011101001",
    "1111001010101101",
    "1111000100101100",
    "1111000001110000",
    "1111000001110100",
    "1111000100101111",
    "1111001010001001",
    "1111010001001111",
    "1111011001000001",
    "1111100000011001",
    "1111100110101111",
    "1111101011110100",
    "1111110000000010",
    "1111110100000000",
    "1111111000011001",
    "1111111101101010",
    "1111111100000011",
    "1111110101001010",
    "1111101110001111",
    "1111101000000000",
    "1111100011001011",
    "1111100000001100",
    "1111011111001000",
    "1111011111110110",
    "1111100001111011",
    "1111100101001000",
    "1111101001100011",
    "1111101111110011",
    "1111111000100100",
    "1111111011110100",
    "1111101101111111",
    "1111011111010110",
    "1111010001110100",
    "1111000111001001",
    "1111000000010111",
    "1110111101010100",
    "1110111100111000",
    "1110111101011011",
    "1110111101101001",
    "1110111101000101",
    "1110111100000111",
    "1110111011101010",
    "1110111100111010",
    "1111000000110110",
    "1111001000001011",
    "1111010011000101",
    "1111100001010000",
    "1111110001111101",
    "1111111100001010",
    "1111101010101011",
    "1111011010111010",
    "1111001101110011",
    "1111000011101110",
    "1110111100100000",
    "1110110111100111",
    "1110110100100010",
    "1110110010111001",
    "1110110010011101",
    "1110110011000001",
    "1110110100001101",
    "1110110101011111",
    "1110110110010010",
    "1110110110000100",
    "1110110100100101",
    "1110110001110110",
    "1110101110010001",
    "1110101010011000",
    "1110100110110110",
    "1110100100001000",
    "1110100010100100",
    "1110100010010101",
    "1110100011100010",
    "1110100110010011",
    "1110101010101101",
    "1110110000110001",
    "1110111000011000",
    "1111000001010100",
    "1111001011011001",
    "1111010110010010",
    "1111100001011001",
    "1111101011111010",
    "1111110101000101",
    "1111111100011111",
    "1111111101110001",
    "1111111000111001",
    "1111110011011101",
    "1111101100000010",
    "1111100001111000",
    "1111010101010000",
    "1111000111010101",
    "1110111001110111",
    "1110101110101000",
    "1110100110110100",
    "1110100010110001",
    "1110100001110100",
    "1110100010111000",
    "1110100100101010",
    "1110100110010110",
    "1110100111100011",
    "1110101000010011",
    "1110101000101000",
    "1110101000101101",
    "1110101000011000",
    "1110100111011111",
    "1110100110000000",
    "1110100011111001",
    "1110100001010111",
    "1110011110110001",
    "1110011100011110",
    "1110011010110100",
    "1110011001111111",
    "1110011010010001",
    "1110011011101101",
    "1110011110010100",
    "1110100010000110",
    "1110100111001110",
    "1110101110101001",
    "1110111001101111",
    "1111001001100011",
    "1111011101110010",
    "1111110100100011",
    "1111110101001011",
    "1111100010111011",
    "1111010111011011",
    "1111010011111000",
    "1111010111011011",
    "1111011111110011",
    "1111101010010110",
    "1111110100110100",
    "1111111101111100",
    "1111111010101111",
    "1111110101010101",
    "1111110001101100",
    "1111101111110101",
    "1111101111110010",
    "1111110001011011",
    "1111110100010010",
    "1111110111100011",
    "1111111010010001",
    "1111111011101101",
    "1111111011101101",
    "1111111010101100",
    "1111111001011110",
    "1111111000101100",
    "1111111000101101",
    "1111111001100010",
    "1111111010110110",
    "1111111100000111",
    "1111111100110111",
    "1111111100110101",
    "1111111100000111",
    "1111111011001001",
    "1111111010100110",
    "1111111011001011",
    "1111111101011011",
    "1111111110010011",
    "1111111000000111",
    "1111110000010011",
    "1111100111011110",
    "1111011110010111",
    "1111010101110110",
    "1111001110101000",
    "1111001001001110",
    "1111000101100101",
    "1111000011010011",
    "1111000001110000",
    "1111000000100100",
    "1110111111101011",
    "1110111111010010",
    "1110111111101100",
    "1111000000110101",
    "1111000010010010",
    "1111000011010111",
    "1111000011011000",
    "1111000001110110",
    "1110111110111000",
    "1110111011000111",
    "1110110111011111",
    "1110110100110110",
    "1110110011101001",
    "1110110011101111",
    "1110110100100101",
    "1110110101011011",
    "1110110101101001",
    "1110110100111100",
    "1110110011100110",
    "1110110010000011",
    "1110110000111101",
    "1110110000101100",
    "1110110001100001",
    "1110110011010000",
    "1110110101101010",
    "1110111000010101",
    "1110111010110101",
    "1110111100110011",
    "1110111101111010",
    "1110111101110111",
    "1110111100101000",
    "1110111010011001",
    "1110110111110010",
    "1110110101101100",
    "1110110101000011",
    "1110110110101000",
    "1110111010101111",
    "1111000001000011",
    "1111001000110010",
    "1111010000110110",
    "1111011000010011",
    "1111011110010111",
    "1111100010110110",
    "1111100101110110",
    "1111100111110101",
    "1111101001010110",
    "1111101010110011",
    "1111101100011011",
    "1111101110010000",
    "1111101111111111",
    "1111110001001111",
    "1111110001101000",
    "1111110000111100",
    "1111101111001110",
    "1111101100101110",
    "1111101001110100",
    "1111100110111011",
    "1111100100011000",
    "1111100010010100",
    "1111100000100110",
    "1111011110111101",
    "1111011101001110",
    "1111011011001110",
    "1111011000111100",
    "1111010110100010",
    "1111010100000110",
    "1111010010000010",
    "1111010000100111",
    "1111010000010100",
    "1111010001010010",
    "1111010011100100",
    "1111010110111100",
    "1111011011001001",
    "1111011111110001",
    "1111100100011111",
    "1111101001000001",
    "1111101101001110",
    "1111110001000110",
    "1111110100101110",
    "1111111000001011",
    "1111111011100000",
    "1111111110101011",
    "1111111110011001",
    "1111111100000000",
    "1111111010001101",
    "1111111000111001",
    "1111110111101110",
    "1111110110010001",
    "1111110100011001",
    "1111110010010101",
    "1111110000100011",
    "1111101111101010",
    "1111110000010010",
    "1111110010101111",
    "1111110111000101",
    "1111111100111001",
    "1111111100100010",
    "1111110110001100",
    "1111110000111101",
    "1111101101100010",
    "1111101100010100",
    "1111101101001111",
    "1111101111111101",
    "1111110011111001",
    "1111111000011000",
    "1111111100110010",
    "1111111111011010",
    "1111111100101101",
    "1111111011010110",
    "1111111011010000",
    "1111111100000001",
    "1111111100111111",
    "1111111101100001",
    "1111111101000111",
    "1111111011011100",
    "1111111000100000",
    "1111110100011110",
    "1111101111100100",
    "1111101010000011",
    "1111100100000101",
    "1111011101111010",
    "1111011000001000",
    "1111010011010111",
    "1111010000010101",
    "1111001111011110",
    "1111010000100110",
    "1111010011001101",
    "1111010110011011",
    "1111011001011101",
    "1111011011110010",
    "1111011101001110",
    "1111011101111010",
    "1111011110000101",
    "1111011110000101",
    "1111011110010100",
    "1111011111010111",
    "1111100001111011",
    "1111100110011111",
    "1111101101001011",
    "1111110101100001",
    "1111111110100011",
    "1111111000111001",
    "1111110010000011",
    "1111101101101001",
    "1111101011111001",
    "1111101100100011",
    "1111101111010000",
    "1111110011100111",
    "1111111001011111",
    "1111111111001001",
    "1111110110100010",
    "1111101100111111",
    "1111100011001010",
    "1111011001110111",
    "1111010010000110",
    "1111001100101110",
    "1111001010010001",
    "1111001010101000",
    "1111001101000100",
    "1111010000000111",
    "1111010010000000",
    "1111010001000011",
    "1111001100010011",
    "1111000011101111",
    "1110111000011011",
    "1110101011111100",
    "1110011111111111",
    "1110010101111100",
    "1110001110100100",
    "1110001010001001",
    "1110001000011010",
    "1110001001000111",
    "1110001100100000",
    "1110010011001011",
    "1110011101111101",
    "1110101100111000",
    "1110111110111010",
    "1111010001110000",
    "1111100010100100",
    "1111101110110011",
    "1111110100110101",
    "1111110100100110",
    "1111101111001111",
    "1111100110110001",
    "1111011101010100",
    "1111010100100101",
    "1111001101101011",
    "1111001001000001",
    "1111000110110010",
    "1111000111000011",
    "1111001001110000",
    "1111001110101110",
    "1111010101010010",
    "1111011100011100",
    "1111100011000101",
    "1111101000000100",
    "1111101010110110",
    "1111101011100100",
    "1111101010111001",
    "1111101001100111",
    "1111101000000010",
    "1111100110001000",
    "1111100011101110",
    "1111100001000010",
    "1111011110101001",
    "1111011101011001",
    "1111011101110010",
    "1111011111101001",
    "1111100010000000",
    "1111100011011010",
    "1111100010011111",
    "1111011110101001",
    "1111011000100010",
    "1111010001110001",
    "1111001100010111",
    "1111001001110100",
    "1111001010101011",
    "1111001110100100",
    "1111010100100000",
    "1111011011100001",
    "1111100011000001",
    "1111101010110110",
    "1111110011001010",
    "1111111100000101",
    "1111111010100110",
    "1111110001101001",
    "1111101001111011",
    "1111100100010010",
    "1111100001010010",
    "1111100001000111",
    "1111100011010011",
    "1111100111001010",
    "1111101011111010",
    "1111110001001001",
    "1111110110111000",
    "1111111101010110",
    "1111111011011001",
    "1111110011111000",
    "1111101101000101",
    "1111101000001000",
    "1111100101110111",
    "1111100110011101",
    "1111101001001111",
    "1111101101000001",
    "1111110000011100",
    "1111110010101010",
    "1111110011100001",
    "1111110011100101",
    "1111110011101101",
    "1111110100110000",
    "1111110111001100",
    "1111111011000010",
    "1111111111111100",
    "1111111010011101",
    "1111110100011101",
    "1111101101111011",
    "1111100110100111",
    "1111011110011011",
    "1111010101101010",
    "1111001101001001",
    "1111000101101110",
    "1111000000000010",
    "1110111100001100",
    "1110111001110010",
    "1110111000000100",
    "1110110110011010",
    "1110110100011000",
    "1110110010000010",
    "1110101111101011",
    "1110101101101000",
    "1110101100000101",
    "1110101011000001",
    "1110101010010011",
    "1110101001111001",
    "1110101001110111",
    "1110101010011000",
    "1110101011100000",
    "1110101101000000",
    "1110101110100110",
    "1110101111101011",
    "1110101111110110",
    "1110101110111000",
    "1110101101000000",
    "1110101010101011",
    "1110101000011101",
    "1110100110101100",
    "1110100101100111",
    "1110100101010000",
    "1110100101101001",
    "1110100110110010",
    "1110101000110010",
    "1110101011101011",
    "1110101111010111",
    "1110110011101010",
    "1110111000010000",
    "1110111100110010",
    "1111000001101110",
    "1111001001001001",
    "1111010101110100",
    "1111101001110011",
    "1111111011000011",
    "1111011011111100",
    "1110111101111000",
    "1110100110010011",
    "1110011001001011",
    "1110010111001001",
    "1110011101101000",
    "1110100111111110",
    "1110110001011110",
    "1110110111000001",
    "1110110111110101",
    "1110110100111110",
    "1110110000010111",
    "1110101011111101",
    "1110101000110010",
    "1110100110111111",
    "1110100110000011",
    "1110100101010101",
    "1110100100101001",
    "1110100100001110",
    "1110100100011101",
    "1110100101011101",
    "1110100110111110",
    "1110101000100011",
    "1110101010001100",
    "1110101100010110",
    "1110110000010111",
    "1110110111111111",
    "1111000100010000",
    "1111010100110110",
    "1111100111110101",
    "1111111010000110",
    "1111110111011011",
    "1111101111001000",
    "1111101101011110",
    "1111110001001100",
    "1111111000000010",
    "1111111111101100",
    "1111111001010101",
    "1111110011100010",
    "1111101110101000",
    "1111101010001100",
    "1111100101111100",
    "1111100010000101",
    "1111011111000111",
    "1111011101100001",
    "1111011101101000",
    "1111011111011111",
    "1111100010101111",
    "1111100110110001",
    "1111101010110110",
    "1111101110010001",
    "1111110000011110",
    "1111110001000111",
    "1111110000001111",
    "1111101110001111",
    "1111101011110111",
    "1111101001111100",
    "1111101001000010",
    "1111101001010011",
    "1111101010011001",
    "1111101011110011",
    "1111101100111110",
    "1111101101101101",
    "1111101110001100",
    "1111101111000101",
    "1111110001010100",
    "1111110101101100",
    "1111111100011110",
    "1111111010101111",
    "1111110001001010",
    "1111101000010000",
    "1111100001010101",
    "1111011101010001",
    "1111011100000101",
    "1111011101010100",
    "1111100000001111",
    "1111100100000011",
    "1111101000000001",
    "1111101011010110",
    "1111101101000111",
    "1111101100011011",
    "1111101000100101",
    "1111100001010100",
    "1111010111000001",
    "1111001010100101",
    "1110111101001111",
    "1110110000010111",
    "1110100100110111",
    "1110011011000111",
    "1110010011000110",
    "1110001100011110",
    "1110000110111001",
    "1110000010001101",
    "1101111110011100",
    "1101111011111101",
    "1101111011000111",
    "1101111100000100",
    "1101111110110110",
    "1110000011001101",
    "1110001000101100",
    "1110001110110101",
    "1110010101010111",
    "1110011100010001",
    "1110100011111000",
    "1110101100101000",
    "1110110110110100",
    "1111000010011001",
    "1111001111000100",
    "1111011100010100",
    "1111101001100110",
    "1111110110010010",
    "1111111110000100",
    "1111110011110100",
    "1111101011000011",
    "1111100011100110",
    "1111011101000100",
    "1111010111000011",
    "1111010001000101",
    "1111001011000111",
    "1111000101010011",
    "1111000000000111",
    "1110111011111101",
    "1110111001001100",
    "1110110111111010",
    "1110111000000110",
    "1110111001101000",
    "1110111100100101",
    "1111000001000011",
    "1111000111011000",
    "1111001111110001",
    "1111011010010011",
    "1111100110101000",
    "1111110100001101",
    "1111111101110000",
    "1111110000010010",
    "1111100100001110",
    "1111011010010110",
    "1111010011001000",
    "1111001110101110",
    "1111001100111100",
    "1111001101001010",
    "1111001110110011",
    "1111010001010000",
    "1111010100000011",
    "1111010110111001",
    "1111011001101010",
    "1111011100010111",
    "1111011111000101",
    "1111100001111011",
    "1111100101000110",
    "1111101000110100",
    "1111101101010001",
    "1111110010011101",
    "1111111000001001",
    "1111111101110010",
    "1111111101010001",
    "1111111001110010",
    "1111111000001100",
    "1111111000101100",
    "1111111011000001",
    "1111111110110000",
    "1111111100011101",
    "1111110110111110",
    "1111110001000000",
    "1111101010111010",
    "1111100101011101",
    "1111100001100110",
    "1111100000001101",
    "1111100001111000",
    "1111100110010011",
    "1111101100101010",
    "1111110011100001",
    "1111111001011001",
    "1111111101000010",
    "1111111101110100",
    "1111111011110100",
    "1111110111101011",
    "1111110010011011",
    "1111101101010011",
    "1111101001011001",
    "1111100111100011",
    "1111101000010100",
    "1111101011111100",
    "1111110010011000",
    "1111111011001101",
    "1111111010010110",
    "1111101111101010",
    "1111100110010011",
    "1111011111111101",
    "1111011101110101",
    "1111100000011100",
    "1111100111001100",
    "1111110000101000",
    "1111111010110010",
    "1111111100001011",
    "1111110101100111",
    "1111110010000100",
    "1111110001011011",
    "1111110011011001",
    "1111110111101001",
    "1111111101111001",
    "1111111010001111",
    "1111110001101100",
    "1111101001110100",
    "1111100100010000",
    "1111100010010101",
    "1111100100101100",
    "1111101010111110",
    "1111110011111010",
    "1111111101110011",
    "1111111001000001",
    "1111110001111101",
    "1111101101110001",
    "1111101100110010",
    "1111101111000101",
    "1111110100101000",
    "1111111101001010",
    "1111110111110101",
    "1111101011100011",
    "1111011111101001",
    "1111010110000011",
    "1111010000101110",
    "1111010000111101",
    "1111010111000001",
    "1111100001111110",
    "1111101111110000",
    "1111111101111101",
    "1111110101100010",
    "1111101100001110",
    "1111100110100110",
    "1111100100011100",
    "1111100101001011",
    "1111101000011010",
    "1111101110001001",
    "1111110110100100",
    "1111111110011100",
    "1111110001111001",
    "1111100101100010",
    "1111011011100110",
    "1111010110010101",
    "1111010111001001",
    "1111011110001010",
    "1111101010000000",
    "1111111000010101",
    "1111111001011111",
    "1111101101110100",
    "1111100101111001",
    "1111100010000110",
    "1111100010000000",
    "1111100100110110",
    "1111101001111011",
    "1111110000101111",
    "1111111000111100",
    "1111111101110010",
    "1111110100000110",
    "1111101010100111",
    "1111100001111000",
    "1111011010010011",
    "1111010100000011",
    "1111001111010010",
    "1111001100000001",
    "1111001010001011",
    "1111001001101010",
    "1111001010011001",
    "1111001100010111",
    "1111001111011110",
    "1111010011011111",
    "1111011000010000",
    "1111011101100011",
    "1111100011010000",
    "1111101001001111",
    "1111101111011000",
    "1111110101011001",
    "1111111010110101",
    "1111111111000011",
    "1111111110101010",
    "1111111111000010",
    "1111111101101010",
    "1111110111101111",
    "1111101111111001",
    "1111100110111110",
    "1111011101110000",
    "1111010100101100",
    "1111001100001001",
    "1111000100010111",
    "1110111101101101",
    "1110111000110000",
    "1110110110001011",
    "1110110110100000",
    "1110111001111101",
    "1111000000001000",
    "1111001000010001",
    "1111010001101100",
    "1111011011111000",
    "1111100110101000",
    "1111110001101110",
    "1111111100110101",
    "1111111000101000",
    "1111101111100100",
    "1111101000101111",
    "1111100100100101",
    "1111100011000000",
    "1111100011011101",
    "1111100101001011",
    "1111100111011110",
    "1111101010000000",
    "1111101100110111",
    "1111110000011011",
    "1111110101000110",
    "1111111011001111",
    "1111111101001101",
    "1111110100110100",
    "1111101100011101",
    "1111100101000011",
    "1111011111010010",
    "1111011011011101",
    "1111011001010101",
    "1111011000010001",
    "1111010111100010",
    "1111010110010110",
    "1111010100010000",
    "1111010001000011",
    "1111001100110101",
    "1111000111110001",
    "1111000010001101",
    "1110111100101010",
    "1110110111101111",
    "1110110100011010",
    "1110110011101110",
    "1110110110110100",
    "1110111110101110",
    "1111001011110111",
    "1111011101101001",
    "1111110010011100",
    "1111111000000100",
    "1111100100010011",
    "1111010011111011",
    "1111000111101101",
    "1110111111011110",
    "1110111010011001",
    "1110110111011011",
    "1110110101101111",
    "1110110100110100",
    "1110110100011111",
    "1110110100101001",
    "1110110101000110",
    "1110110101101010",
    "1110110110001011",
    "1110110110011011",
    "1110110110011010",
    "1110110110001001",
    "1110110101101110",
    "1110110101001011",
    "1110110100100010",
    "1110110011110001",
    "1110110010111001",
    "1110110010000011",
    "1110110001100110",
    "1110110001111110",
    "1110110011011111",
    "1110110110010011",
    "1110111010010001",
    "1110111111001100",
    "1111000100101010",
    "1111001010010011",
    "1111001111101100",
    "1111010100011111",
    "1111011000011011",
    "1111011011110000",
    "1111011111100011",
    "1111100101100000",
    "1111101111010000",
    "1111111101101110",
    "1111101111101010",
    "1111011010111101",
    "1111000111001011",
    "1110110111011010",
    "1110101101101011",
    "1110101010001100",
    "1110101011100001",
    "1110101111001101",
    "1110110010101011",
    "1110110100000101",
    "1110110010110011",
    "1110101111001111",
    "1110101010011101",
    "1110100101011101",
    "1110100000111001",
    "1110011101001001",
    "1110011010000001",
    "1110010111011111",
    "1110010101011101",
    "1110010100000011",
    "1110010011011000",
    "1110010011011010",
    "1110010100000011",
    "1110010101000110",
    "1110010110010110",
    "1110010111101100",
    "1110011001000111",
    "1110011010110010",
    "1110011101001001",
    "1110100000111110",
    "1110100111100010",
    "1110110001110110",
    "1111000000000111",
    "1111010001001101",
    "1111100010111000",
    "1111110010010001",
    "1111111100111101",
    "1111111110010101",
    "1111111111010000",
    "1111111100000111",
    "1111110110011010",
    "1111110001110110",
    "1111101111101010",
    "1111101111110101",
    "1111110001011111",
    "1111110011100001",
    "1111110101000101",
    "1111110101111010",
    "1111110110001100",
    "1111110110010011",
    "1111110110011011",
    "1111110110100011",
    "1111110110011100",
    "1111110101111000",
    "1111110100111110",
    "1111110011111101",
    "1111110011001010",
    "1111110010101111",
    "1111110010100110",
    "1111110010100010",
    "1111110010010101",
    "1111110001111110",
    "1111110001101000",
    "1111110001100100",
    "1111110010001100",
    "1111110011111001",
    "1111110110111110",
    "1111111011101001",
    "1111111101111110",
    "1111110110000111",
    "1111101101001000",
    "1111100011101010",
    "1111011010011110",
    "1111010010001101",
    "1111001011011011",
    "1111000110011101",
    "1111000011011000",
    "1111000010001011",
    "1111000010101001",
    "1111000100010111",
    "1111000110110110",
    "1111001001011001",
    "1111001011010110",
    "1111001100001100",
    "1111001011101010",
    "1111001001110111",
    "1111000111010011",
    "1111000100011111",
    "1111000001111101",
    "1111000000000000",
    "1110111110110001",
    "1110111110001100",
    "1110111101111111",
    "1110111101110011",
    "1110111101010001",
    "1110111100000010",
    "1110111001111010",
    "1110110111000110",
    "1110110011111110",
    "1110110001001000",
    "1110101111001100",
    "1110101110011100",
    "1110101111000010",
    "1110110000101100",
    "1110110011000011",
    "1110110101100010",
    "1110110111101100",
    "1110111001000100",
    "1110111001011001",
    "1110111000110100",
    "1110110111101010",
    "1110110110100100",
    "1110110110000000",
    "1110110110010010",
    "1110110111010110",
    "1110111001000111",
    "1110111011101010",
    "1110111111001010",
    "1111000100000101",
    "1111001010110000",
    "1111010011000001",
    "1111011100001010",
    "1111100101000001",
    "1111101100010011",
    "1111110001010000",
    "1111110011101111",
    "1111110100001101",
    "1111110011011111",
    "1111110010011100",
    "1111110001101100",
    "1111110001100001",
    "1111110001111001",
    "1111110010100110",
    "1111110011011110",
    "1111110100010011",
    "1111110100101111",
    "1111110100010001",
    "1111110010010001",
    "1111101110001110",
    "1111100111111100",
    "1111011111101000",
    "1111010110000110",
    "1111001100100110",
    "1111000100011111",
    "1110111110111011",
    "1110111100100110",
    "1110111101100001",
    "1111000001001111",
    "1111000111000110",
    "1111001110011001",
    "1111010110100000",
    "1111011110110101",
    "1111100110101000",
    "1111101101010010",
    "1111110010000100",
    "1111110100010110",
    "1111110011111100",
    "1111110001010000",
    "1111101101010110",
    "1111101001101001",
    "1111100111101100",
    "1111101000101101",
    "1111101101001110",
    "1111110100111100",
    "1111111110101110",
    "1111110111000011",
    "1111101110001011",
    "1111100111111001",
    "1111100100110111",
    "1111100101010000",
    "1111101000110111",
    "1111101111011001",
    "1111111000011001",
    "1111111100110110",
    "1111110001100000",
    "1111100110111011",
    "1111011110100110",
    "1111011001110111",
    "1111011001011101",
    "1111011101010100",
    "1111100100100111",
    "1111101110000101",
    "1111111000000111",
    "1111111110110111",
    "1111111000010010",
    "1111110100111111",
    "1111110101010010",
    "1111111000110101",
    "1111111110101001",
    "1111111010100001",
    "1111110100001010",
    "1111101111100001",
    "1111101101011101",
    "1111101110011110",
    "1111110010100011",
    "1111111001011111",
    "1111111101001110",
    "1111110010011010",
    "1111100111000101",
    "1111011100100000",
    "1111010011111011",
    "1111001110010111",
    "1111001100011001",
    "1111001101111101",
    "1111010010011111",
    "1111011000111110",
    "1111100000001101",
    "1111100111000110",
    "1111101100101101",
    "1111110000011000",
    "1111110001110010",
    "1111110000111100",
    "1111101110001000",
    "1111101001111010",
    "1111100101001000",
    "1111100000110011",
    "1111011110000101",
    "1111011110000111",
    "1111100001100001",
    "1111101000011001",
    "1111110010000010",
    "1111111101001110",
    "1111110111011011",
    "1111101101010100",
    "1111100101010111",
    "1111011111111101",
    "1111011101000101",
    "1111011100100000",
    "1111011101110111",
    "1111100001000101",
    "1111100110001110",
    "1111101101011100",
    "1111110110110010",
    "1111111101111100",
    "1111110001011111",
    "1111100100101010",
    "1111011000011010",
    "1111001101100001",
    "1111000100100101",
    "1110111101111011",
    "1110111001100101",
    "1110110111010001",
    "1110110110101000",
    "1110110111000011",
    "1110110111110101",
    "1110111000010110",
    "1110111000001110",
    "1110110111010110",
    "1110110101111110",
    "1110110100100010",
    "1110110011011010",
    "1110110010111000",
    "1110110010111110",
    "1110110011100010",
    "1110110100010011",
    "1110110101000110",
    "1110110101110111",
    "1110110110100101",
    "1110110111001101",
    "1110110111101100",
    "1110110111111001",
    "1110110111111010",
    "1110111000000100",
    "1110111000111001",
    "1110111010111000",
    "1110111110100100",
    "1111000100001000",
    "1111001011011001",
    "1111010011111011",
    "1111011101000100",
    "1111100110001011",
    "1111101110011111",
    "1111110101010110",
    "1111111010000101",
    "1111111100010011",
    "1111111011111101",
    "1111111001010111",
    "1111110101000101",
    "1111101111110010",
    "1111101010000011",
    "1111100100001101",
    "1111011110011001",
    "1111011000100011",
    "1111010010101111",
    "1111001101001001",
    "1111001000000110",
    "1111000100000001",
    "1111000001010000",
    "1110111111111111",
    "1111000000001101",
    "1111000001111101",
    "1111000101010000",
    "1111001010001100",
    "1111010000110110",
    "1111011001001011",
    "1111100010111110",
    "1111101101110011",
    "1111111000110111",
    "1111111100110000",
    "1111110100000100",
    "1111101101110010",
    "1111101010001111",
    "1111101001010110",
    "1111101010100100",
    "1111101101001001",
    "1111110000010010",
    "1111110011011001",
    "1111110110001010",
    "1111111000100011",
    "1111111010101100",
    "1111111100110011",
    "1111111111000000",
    "1111111110100011",
    "1111111011111110",
    "1111111001010111",
    "1111110110111100",
    "1111110100111010",
    "1111110011011000",
    "1111110010010101",
    "1111110001100011",
    "1111110000101011",
    "1111101111010100",
    "1111101101001110",
    "1111101010011010",
    "1111100111001011",
    "1111100100000000",
    "1111100001011110",
    "1111100000000011",
    "1111100000001000",
    "1111100010000010",
    "1111100101111100",
    "1111101100010001",
    "1111110101010110",
    "1111111110100001",
    "1111101111100010",
    "1111011110011111",
    "1111001101000010",
    "1110111101001110",
    "1110110000110110",
    "1110101000111111",
    "1110100101101010",
    "1110100101111100",
    "1110101000010110",
    "1110101011100000",
    "1110101110010111",
    "1110110000101110",
    "1110110010100111",
    "1110110100010111",
    "1110110110000000",
    "1110110111011010",
    "1110111000010001",
    "1110111000010001",
    "1110110111010001",
    "1110110101011000",
    "1110110010111101",
    "1110110000011001",
    "1110101110000000",
    "1110101100000010",
    "1110101010100000",
    "1110101001011011",
    "1110101000111010",
    "1110101001001011",
    "1110101010010110",
    "1110101100100000",
    "1110101111011110",
    "1110110010111101",
    "1110110110100100",
    "1110111001110101",
    "1110111100010110",
    "1110111101110101",
    "1110111110001101",
    "1110111101100110",
    "1110111100001111",
    "1110111010100011",
    "1110111001000100",
    "1110111000010110",
    "1110111001101101",
    "1110111111110101",
    "1111001101101101",
    "1111100100111100",
    "1111111011011011",
    "1111010111100000",
    "1110110101000011",
    "1110011001111001",
    "1110001001111111",
    "1110000101111100",
    "1110001010111101",
    "1110010100011100",
    "1110011101110000",
    "1110100100000001",
    "1110100110011111",
    "1110100101111001",
    "1110100011111001",
    "1110100010000011",
    "1110100001000011",
    "1110100000110011",
    "1110100000111101",
    "1110100001000011",
    "1110100001001010",
    "1110100001100100",
    "1110100010101001",
    "1110100100010101",
    "1110100110001000",
    "1110100111100101",
    "1110101000101000",
    "1110101001101000",
    "1110101011010110",
    "1110101110111111",
    "1110110101101010",
    "1110111111110000",
    "1111001100101110",
    "1111011011000110",
    "1111101000110001",
    "1111110011111010",
    "1111111011001000",
    "1111111101110110",
    "1111111100011101",
    "1111110111110110",
    "1111110001001110",
    "1111101001110010",
    "1111100010101001",
    "1111011100111100",
    "1111011001100111",
    "1111011000111111",
    "1111011010111000",
    "1111011110011100",
    "1111100010100001",
    "1111100110001000",
    "1111101000100010",
    "1111101001100000",
    "1111101001001011",
    "1111100111111011",
    "1111100110001110",
    "1111100100011101",
    "1111100010110011",
    "1111100001011001",
    "1111100000100011",
    "1111100000110000",
    "1111100010011100",
    "1111100101101111",
    "1111101010010010",
    "1111101111011101",
    "1111110100100011",
    "1111111001000100",
    "1111111100110111",
    "1111111111101001",
    "1111111011111110",
    "1111110111011100",
    "1111110001110010",
    "1111101011001100",
    "1111100100011000",
    "1111011110011001",
    "1111011010010110",
    "1111011001000110",
    "1111011010110100",
    "1111011111001010",
    "1111100101001101",
    "1111101011111010",
    "1111110010010001",
    "1111110111011011",
    "1111111010101100",
    "1111111011011010",
    "1111111000110110",
    "1111110010011010",
    "1111100111110010",
    "1111011001010011",
    "1111001000001011",
    "1110110110010110",
    "1110100101111100",
    "1110011000101010",
    "1110001111001111",
    "1110001001011101",
    "1110000110001011",
    "1110000100000000",
    "1110000001110100",
    "1101111111000111",
    "1101111100000111",
    "1101111001011101",
    "1101110111110010",
    "1101110111101100",
    "1101111001001110",
    "1101111100001111",
    "1110000000100001",
    "1110000101110100",
    "1110001100010011",
    "1110010100010011",
    "1110011110001100",
    "1110101001110101",
    "1110110110101101",
    "1111000011110110",
    "1111010000001111",
    "1111011011001100",
    "1111100100100100",
    "1111101100110101",
    "1111110100110001",
    "1111111101001100",
    "1111111001011011",
    "1111101111001011",
    "1111100100011000",
    "1111011001101010",
    "1111001111011111",
    "1111000110010011",
    "1110111110010111",
    "1110110111111010",
    "1110110011001011",
    "1110110000011110",
    "1110110000001111",
    "1110110011000001",
    "1110111001010110",
    "1111000011011111",
    "1111010001010100",
    "1111100001111101",
    "1111110011111101",
    "1111111010100001",
    "1111101011011100",
    "1111100000001101",
    "1111011001011101",
    "1111010110110100",
    "1111010111010000",
    "1111011001011110",
    "1111011100001010",
    "1111011110010001",
    "1111011111001010",
    "1111011110101000",
    "1111011100111100",
    "1111011010100011",
    "1111011000001001",
    "1111010110011011",
    "1111010110001011",
    "1111010111111111",
    "1111011100001111",
    "1111100010111101",
    "1111101011101010",
    "1111110101100000",
    "1111111111010001",
    "1111111000010010",
    "1111110010011000",
    "1111101111110011",
    "1111110000111101",
    "1111110101101111",
    "1111111101101001",
    "1111111000010101",
    "1111101101100111",
    "1111100011101111",
    "1111011100001110",
    "1111011000001001",
    "1111010111111110",
    "1111011011011011",
    "1111100001100110",
    "1111101001001100",
    "1111110000111001",
    "1111110111100110",
    "1111111100011101",
    "1111111110111110",
    "1111111110110110",
    "1111111100000011",
    "1111110110111000",
    "1111110000000111",
    "1111101000111110",
    "1111100010111011",
    "1111011111010111",
    "1111011111001101",
    "1111100010110001",
    "1111101001110110",
    "1111110011110000",
    "1111111111100010",
    "1111110011110110",
    "1111100111100100",
    "1111011100110010",
    "1111010100100101",
    "1111001111111111",
    "1111001111101110",
    "1111010100000110",
    "1111011100111000",
    "1111101001000011",
    "1111110110111101",
    "1111111011010101",
    "1111101111110110",
    "1111101000000001",
    "1111100100100010",
    "1111100101010011",
    "1111101001101000",
    "1111110000100101",
    "1111111001001110",
    "1111111101000110",
    "1111110011000110",
    "1111101001010111",
    "1111100000101110",
    "1111011010000111",
    "1111010110100100",
    "1111010110101111",
    "1111011010101101",
    "1111100001111000",
    "1111101010111100",
    "1111110100011100",
    "1111111100111111",
    "1111111100001111",
    "1111110111110000",
    "1111110101011101",
    "1111110101000000",
    "1111110101111010",
    "1111110111101101",
    "1111111001111111",
    "1111111100011100",
    "1111111110111000",
    "1111111110101110",
    "1111111100100000",
    "1111111010011010",
    "1111111000011111",
    "1111110110110001",
    "1111110101010000",
    "1111110011111011",
    "1111110010110010",
    "1111110001110101",
    "1111110001001111",
    "1111110001010100",
    "1111110010100000",
    "1111110101010011",
    "1111111010000100",
    "1111111111010010",
    "1111110111011010",
    "1111101111010000",
    "1111100111111111",
    "1111100010100111",
    "1111011111111011",
    "1111100000001100",
    "1111100011001101",
    "1111101000100010",
    "1111101111011110",
    "1111110111010011",
    "1111111111011000",
    "1111111000101110",
    "1111110001001100",
    "1111101001110101",
    "1111100010010000",
    "1111011010001110",
    "1111010001110110",
    "1111001001110100",
    "1111000011000110",
    "1110111110110101",
    "1110111101101101",
    "1111000000000010",
    "1111000101100111",
    "1111001101101011",
    "1111010111001110",
    "1111100001001101",
    "1111101010100111",
    "1111110010100111",
    "1111111000100100",
    "1111111100001001",
    "1111111101011100",
    "1111111100110110",
    "1111111010111101",
    "1111111000001101",
    "1111110100110011",
    "1111110000101000",
    "1111101011010111",
    "1111100100101111",
    "1111011100101101",
    "1111010011100100",
    "1111001001111100",
    "1111000000110001",
    "1110111000111001",
    "1110110011000101",
    "1110101111110000",
    "1110101111000101",
    "1110110000111110",
    "1110110101000011",
    "1110111010110101",
    "1111000001111011",
    "1111001001111101",
    "1111010010110001",
    "1111011100001010",
    "1111100101110100",
    "1111101111001100",
    "1111110111011111",
    "1111111101111010",
    "1111111101111101",
    "1111111100001101",
    "1111111100010000",
    "1111111101001110",
    "1111111110000111",
    "1111111110001011",
    "1111111101000100",
    "1111111010110110",
    "1111111000000000",
    "1111110101001100",
    "1111110011001000",
    "1111110010010111",
    "1111110011001111",
    "1111110101111000",
    "1111111010010001",
    "1111111111101011",
    "1111111000001100",
    "1111101111100000",
    "1111100101111110",
    "1111011100000111",
    "1111010010011101",
    "1111001001100011",
    "1111000001101110",
    "1110111011000100",
    "1110110101100000",
    "1110110001000011",
    "1110101101101110",
    "1110101011111100",
    "1110101100001100",
    "1110101111000111",
    "1110110101001000",
    "1110111110001101",
    "1111001010000010",
    "1111010111110111",
    "1111100110101111",
    "1111110101100100",
    "1111111100100111",
    "1111110000101111",
    "1111100111001101",
    "1111011111111111",
    "1111011010100011",
    "1111010110000110",
    "1111010001110011",
    "1111001101000111",
    "1111000111111010",
    "1111000010011100",
    "1110111101001010",
    "1110111000011101",
    "1110110100100010",
    "1110110001011010",
    "1110101111000010",
    "1110101101010100",
    "1110101100001111",
    "1110101011111000",
    "1110101100010111",
    "1110101101101011",
    "1110101111101100",
    "1110110010010010",
    "1110110101001001",
    "1110110111111111",
    "1110111010101011",
    "1110111101001001",
    "1110111111011010",
    "1111000001100111",
    "1111000011110110",
    "1111000110001000",
    "1111001000011010",
    "1111001010100011",
    "1111001100011001",
    "1111001101101110",
    "1111001110011111",
    "1111001110101001",
    "1111001110010100",
    "1111001110101000",
    "1111010010000000",
    "1111011011010001",
    "1111101100001101",
    "1111111011110010",
    "1111011111111011",
    "1111000100111001",
    "1110101111011111",
    "1110100011000110",
    "1110100000000101",
    "1110100100000000",
    "1110101010111100",
    "1110110001000011",
    "1110110100000001",
    "1110110011011000",
    "1110110000000010",
    "1110101011011101",
    "1110100111000011",
    "1110100011011000",
    "1110100000011110",
    "1110011101111011",
    "1110011011011011",
    "1110011001000111",
    "1110010111010110",
    "1110010110011011",
    "1110010110010011",
    "1110010110100010",
    "1110010110101111",
    "1110010110110100",
    "1110010111000001",
    "1110010111101100",
    "1110011001010011",
    "1110011100001010",
    "1110100000011111",
    "1110100110011101",
    "1110101110010010",
    "1110111000001011",
    "1111000100001000",
    "1111010001101011",
    "1111011111101100",
    "1111101100100100",
    "1111110110100101",
    "1111111100011001",
    "1111111101101000",
    "1111111010111110",
    "1111110110001000",
    "1111110001001111",
    "1111101110000100",
    "1111101101100001",
    "1111101111100000",
    "1111110011000110",
    "1111110111000110",
    "1111111010010111",
    "1111111100001000",
    "1111111100000101",
    "1111111010010101",
    "1111110111010010",
    "1111110011100010",
    "1111101111101001",
    "1111101100000110",
    "1111101001010111",
    "1111100111110111",
    "1111100111110101",
    "1111101001010101",
    "1111101100001100",
    "1111110000000111",
    "1111110100110000",
    "1111111001110000",
    "1111111110110010",
    "1111111100001101",
    "1111110111010010",
    "1111110010001111",
    "1111101100111010",
    "1111100111001101",
    "1111100001001000",
    "1111011010111000",
    "1111010100101111",
    "1111001111000101",
    "1111001010001111",
    "1111000110011010",
    "1111000011101100",
    "1111000010000011",
    "1111000001010111",
    "1111000001100010",
    "1111000010011010",
    "1111000011111100",
    "1111000110000001",
    "1111001000010110",
    "1111001010100000",
    "1111001011111000",
    "1111001011111111",
    "1111001010100101",
    "1111000111110100",
    "1111000100001010",
    "1111000000001101",
    "1110111100011011",
    "1110111001000010",
    "1110110110000000",
    "1110110011001010",
    "1110110000011110",
    "1110101110000101",
    "1110101100100000",
    "1110101100001010",
    "1110101101011011",
    "1110110000001000",
    "1110110011110100",
    "1110110111100101",
    "1110111010011101",
    "1110111011100011",
    "1110111010011101",
    "1110110111001011",
    "1110110010001010",
    "1110101100000111",
    "1110100110000011",
    "1110100000111001",
    "1110011101101000",
    "1110011100111100",
    "1110011111010001",
    "1110100100101111",
    "1110101101001110",
    "1110111000001000",
    "1111000100100010",
    "1111010001001100",
    "1111011100101101",
    "1111100101110100",
    "1111101011100101",
    "1111101101110000",
    "1111101100110000",
    "1111101001100011",
    "1111100101100000",
    "1111100001111110",
    "1111100000000111",
    "1111100000011111",
    "1111100011010101",
    "1111101000010011",
    "1111101110100101",
    "1111110101000011",
    "1111111010011000",
    "1111111101010000",
    "1111111100101010",
    "1111111000001000",
    "1111101111111011",
    "1111100101000001",
    "1111011001000001",
    "1111001101100011",
    "1111000011111100",
    "1110111101000100",
    "1110111001000100",
    "1110110111110010",
    "1110111000111111",
    "1110111100011100",
    "1111000010000000",
    "1111001001011101",
    "1111010010010101",
    "1111011011110000",
    "1111100100100100",
    "1111101011010101",
    "1111101111000000",
    "1111101111000110",
    "1111101011111111",
    "1111100110110100",
    "1111100001001111",
    "1111011100110111",
    "1111011010111101",
    "1111011100010011",
    "1111100000111000",
    "1111101000010011",
    "1111110001110101",
    "1111111100100110",
    "1111111000011101",
    "1111101110100100",
    "1111100110111001",
    "1111100010100111",
    "1111100010101001",
    "1111100111011010",
    "1111110000100101",
    "1111111100111111",
    "1111110101000111",
    "1111100111110011",
    "1111011100110000",
    "1111010101001101",
    "1111010001110100",
    "1111010010101011",
    "1111010111100010",
    "1111011111111011",
    "1111101011000110",
    "1111110111111011",
    "1111111010111110",
    "1111101111010001",
    "1111100110011100",
    "1111100001011110",
    "1111100000111000",
    "1111100100100100",
    "1111101011110010",
    "1111110101010001",
    "1111111111011100",
    "1111110111010001",
    "1111110000010011",
    "1111101100011110",
    "1111101100000100",
    "1111101110110011",
    "1111110100000001",
    "1111111010111101",
    "1111111100111100",
    "1111110100001010",
    "1111101010111010",
    "1111100001011110",
    "1111011000000100",
    "1111001111001010",
    "1111000111010000",
    "1111000000110110",
    "1110111100011110",
    "1110111010100000",
    "1110111011001110",
    "1110111110101101",
    "1111000100110011",
    "1111001101001010",
    "1111010111010000",
    "1111100010011001",
    "1111101101110011",
    "1111111000110010",
    "1111111101001110",
    "1111110100110010",
    "1111101110001011",
    "1111101001100000",
    "1111100110101111",
    "1111100101101100",
    "1111100110001000",
    "1111100111110010",
    "1111101010011100",
    "1111101101110111",
    "1111110001110100",
    "1111110110000011",
    "1111111010010110",
    "1111111110100100",
    "1111111101011000",
    "1111111001100110",
    "1111110110001000",
    "1111110011000100",
    "1111110000100101",
    "1111101110101101",
    "1111101101010101",
    "1111101100001010",
    "1111101010110010",
    "1111101000101111",
    "1111100101101110",
    "1111100001100010",
    "1111011100010011",
    "1111010110000011",
    "1111001110111011",
    "1111000111000011",
    "1110111110100011",
    "1110110101111001",
    "1110101101100100",
    "1110100110010011",
    "1110100000101001",
    "1110011100110101",
    "1110011010110100",
    "1110011010000111",
    "1110011010000111",
    "1110011010001111",
    "1110011010001111",
    "1110011010010011",
    "1110011011000100",
    "1110011101011100",
    "1110100010001011",
    "1110101001110000",
    "1110110100000001",
    "1111000000010001",
    "1111001101010110",
    "1111011010000111",
    "1111100101100010",
    "1111101110110000",
    "1111110101001011",
    "1111111000100010",
    "1111111000110101",
    "1111110110010111",
    "1111110001110000",
    "1111101011110000",
    "1111100101001011",
    "1111011110101101",
    "1111011000101000",
    "1111010011000000",
    "1111001101100001",
    "1111001000000011",
    "1111000010100100",
    "1110111101011011",
    "1110111001010000",
    "1110110110101010",
    "1110110110001001",
    "1110110111110010",
    "1110111011001111",
    "1110111111111101",
    "1111000101010010",
    "1111001010101000",
    "1111001111110001",
    "1111010100101001",
    "1111011001011000",
    "1111011110000100",
    "1111100010110011",
    "1111100111100010",
    "1111101100010000",
    "1111110001000000",
    "1111110101111010",
    "1111111011001101",
    "1111111111000001",
    "1111111001000001",
    "1111110011001101",
    "1111101110001110",
    "1111101010101111",
    "1111101001001100",
    "1111101001110010",
    "1111101100011110",
    "1111110001000101",
    "1111110111100000",
    "1111111111100010",
    "1111110110111110",
    "1111101100101001",
    "1111100010001101",
    "1111011000101100",
    "1111010001000011",
    "1111001011111111",
    "1111001001101111",
    "1111001001110111",
    "1111001011101011",
    "1111001110010010",
    "1111010001000011",
    "1111010011101001",
    "1111010110000110",
    "1111011000101101",
    "1111011011111101",
    "1111100000001111",
    "1111100101110111",
    "1111101100111101",
    "1111110101100011",
    "1111111111100000",
    "1111110101010100",
    "1111101001010111",
    "1111011101010001",
    "1111010001111001",
    "1111001000001100",
    "1111000000111101",
    "1110111100010110",
    "1110111010001001",
    "1110111001100011",
    "1110111001100101",
    "1110111001011110",
    "1110111000110101",
    "1110110111101101",
    "1110110110100100",
    "1110110101111011",
    "1110110110001101",
    "1110110111100000",
    "1110111001011110",
    "1110111011011110",
    "1110111100101101",
    "1110111100100001",
    "1110111010110100",
    "1110110111110111",
    "1110110100011010",
    "1110110001010010",
    "1110101111001010",
    "1110101110010010",
    "1110101110100110",
    "1110101111101001",
    "1110110000111101",
    "1110110010000011",
    "1110110010101111",
    "1110110011000001",
    "1110110011000000",
    "1110110010110011",
    "1110110010011001",
    "1110110001110001",
    "1110110000111000",
    "1110101111101011",
    "1110101110010001",
    "1110101100111100",
    "1110101011111101",
    "1110101011101111",
    "1110101100101010",
    "1110101111101110",
    "1110110111010001",
    "1111000101111100",
    "1111011101001100",
    "1111111100000111",
    "1111100000111101",
    "1110111111011010",
    "1110100100100101",
    "1110010100001011",
    "1110001110110011",
    "1110010001111000",
    "1110011001000110",
    "1110100000001101",
    "1110100100100111",
    "1110100101101010",
    "1110100100010101",
    "1110100010010101",
    "1110100001001100",
    "1110100001100100",
    "1110100011010000",
    "1110100101100100",
    "1110100111101111",
    "1110101001011101",
    "1110101010110111",
    "1110101100001010",
    "1110101101010111",
    "1110101110001101",
    "1110101110100001",
    "1110101110011100",
    "1110101110011001",
    "1110101111000000",
    "1110110000111000",
    "1110110100101010",
    "1110111010111000",
    "1111000011101010",
    "1111001110101110",
    "1111011011000111",
    "1111100111101011",
    "1111110010111101",
    "1111111011100011",
    "1111111111011100",
    "1111111110011001",
    "1111111111001001",
    "1111111010010001",
    "1111110100001110",
    "1111101110001111",
    "1111101001001101",
    "1111100101100010",
    "1111100011000101",
    "1111100001011010",
    "1111100000010111",
    "1111011111111010",
    "1111100000010010",
    "1111100001101001",
    "1111100011110011",
    "1111100110001110",
    "1111101000011000",
    "1111101001110100",
    "1111101010100001",
    "1111101010101111",
    "1111101011000101",
    "1111101100001111",
    "1111101110101011",
    "1111110010100001",
    "1111110111011101",
    "1111111101000001",
    "1111111101000111",
    "1111110111010010",
    "1111110001011111",
    "1111101011100111",
    "1111100101101001",
    "1111011111101110",
    "1111011010011000",
    "1111010110010110",
    "1111010100100010",
    "1111010101011111",
    "1111011001010101",
    "1111011111100100",
    "1111100111010000",
    "1111101111000101",
    "1111110101110110",
    "1111111010101101",
    "1111111101001101",
    "1111111101001000",
    "1111111010011001",
    "1111110100111111",
    "1111101101000100",
    "1111100011000001",
    "1111010111101100",
    "1111001100000010",
    "1111000001001000",
    "1110110111101100",
    "1110101111111111",
    "1110101001110101",
    "1110100100101100",
    "1110011111110110",
    "1110011010100110",
    "1110010100100111",
    "1110001101101101",
    "1110000110001000",
    "1101111110010111",
    "1101110111001000",
    "1101110001001010",
    "1101101101001001",
    "1101101011100000",
    "1101101100011001",
    "1101101111101110",
    "1101110101010101",
    "1101111100111111",
    "1110000110010110",
    "1110010001000101",
    "1110011100100000",
    "1110100111111010",
    "1110110010101011",
    "1110111100010110",
    "1111000100111100",
    "1111001100111111",
    "1111010101010101",
    "1111011110110101",
    "1111101010000100",
    "1111110111000110",
    "1111111010100011",
    "1111101011111101",
    "1111011110001010",
    "1111010010001000",
    "1111001000010110",
    "1111000001000000",
    "1110111011110011",
    "1110111000010110",
    "1110110110011111",
    "1110110110010110",
    "1110111000101111",
    "1110111110101011",
    "1111001000111010",
    "1111010111010110",
    "1111101000110000",
    "1111111010111110",
    "1111110100100011",
    "1111101000001010",
    "1111100001000101",
    "1111011111010110",
    "1111100001101110",
    "1111100110011010",
    "1111101011011101",
    "1111101111010001",
    "1111110000111100",
    "1111110000001111",
    "1111101101011011",
    "1111101001001100",
    "1111100100010011",
    "1111011111011111",
    "1111011011100000",
    "1111011000111110",
    "1111011000011110",
    "1111011010100000",
    "1111011111001100",
    "1111100110011011",
    "1111101111101011",
    "1111111010001101",
    "1111111011000101",
    "1111110001100001",
    "1111101010011001",
    "1111100110110001",
    "1111100111010100",
    "1111101100000010",
    "1111110100010101",
    "1111111111000110",
    "1111110100111111",
    "1111101001011111",
    "1111011111100100",
    "1111011000001011",
    "1111010011101110",
    "1111010010010010",
    "1111010011100010",
    "1111010110111100",
    "1111011011111000",
    "1111100001110110",
    "1111101000011100",
    "1111101111010111",
    "1111110110010000",
    "1111111100110111",
    "1111111101000000",
    "1111110111101110",
    "1111110011100000",
    "1111110000100011",
    "1111101110111110",
    "1111101110110011",
    "1111101111111100",
    "1111110010001101",
    "1111110101011001",
    "1111111001001000",
    "1111111100111100",
    "1111111111101010",
    "1111111101010101",
    "1111111100011000",
    "1111111100111010",
    "1111111110101100",
    "1111111110101001",
    "1111111011101101",
    "1111111000110111",
    "1111110110010100",
    "1111110100000110",
    "1111110010000011",
    "1111101111111111",
    "1111101101110100",
    "1111101011100101",
    "1111101001011111",
    "1111100111111001",
    "1111100111001010",
    "1111100111100010",
    "1111101001001000",
    "1111101011110111",
    "1111101111100000",
    "1111110011110000",
    "1111111000010100",
    "1111111100110100",
    "1111111111000010",
    "1111111011110000",
    "1111111001101111",
    "1111111001010101",
    "1111111010101110",
    "1111111101111010",
    "1111111101011100",
    "1111111000000000",
    "1111110010011101",
    "1111101101011100",
    "1111101001011001",
    "1111100110011011",
    "1111100100011000",
    "1111100011000110",
    "1111100010100001",
    "1111100010101011",
    "1111100011111000",
    "1111100110011101",
    "1111101010100011",
    "1111101111111100",
    "1111110110001011",
    "1111111100100011",
    "1111111101011110",
    "1111111000011010",
    "1111110100001101",
    "1111110000110001",
    "1111101101110101",
    "1111101011010010",
    "1111101001001111",
    "1111101000000010",
    "1111101000000101",
    "1111101001101110",
    "1111101101001001",
    "1111110010010011",
    "1111111000111110",
    "1111111111001101",
    "1111110110110000",
    "1111101110001001",
    "1111100101110110",
    "1111011110010100",
    "1111011000000011",
    "1111010011011100",
    "1111010000111000",
    "1111010000100011",
    "1111010010010100",
    "1111010101110111",
    "1111011010100110",
    "1111011111110110",
    "1111100101000001",
    "1111101001100111",
    "1111101101010110",
    "1111110000000101",
    "1111110001101101",
    "1111110010001001",
    "1111110001010101",
    "1111101111010110",
    "1111101100011101",
    "1111101001001100",
    "1111100110001000",
    "1111100011110001",
    "1111100010011001",
    "1111100001111001",
    "1111100001111001",
    "1111100001110011",
    "1111100000111000",
    "1111011110101000",
    "1111011010101111",
    "1111010101001011",
    "1111001110010010",
    "1111000110100101",
    "1110111110101110",
    "1110110111010110",
    "1110110001000101",
    "1110101100010110",
    "1110101001100111",
    "1110101001001110",
    "1110101011100101",
    "1110110001000010",
    "1110111001100111",
    "1111000100111100",
    "1111010010010000",
    "1111100000010111",
    "1111101101110111",
    "1111111001100101",
    "1111111101010001",
    "1111110111000001",
    "1111110011010110",
    "1111110001110001",
    "1111110001100110",
    "1111110010011001",
    "1111110011110110",
    "1111110101110111",
    "1111111000011100",
    "1111111011100111",
    "1111111111011010",
    "1111111100001100",
    "1111110111010010",
    "1111110001111100",
    "1111101100011000",
    "1111100110111001",
    "1111100001110001",
    "1111011101010111",
    "1111011001110000",
    "1111010110111001",
    "1111010100010111",
    "1111010001101110",
    "1111001110100110",
    "1111001010110100",
    "1111000110011011",
    "1111000001111000",
    "1110111101101011",
    "1110111010011001",
    "1110111000100011",
    "1110111000100000",
    "1110111010100010",
    "1110111110110011",
    "1111000101011010",
    "1111001110010010",
    "1111011001000110",
    "1111100101001011",
    "1111110001101010",
    "1111111101100000",
    "1111111000000111",
    "1111101111101110",
    "1111101001001111",
    "1111100100000101",
    "1111011111010111",
    "1111011010001110",
    "1111010100001011",
    "1111001101001110",
    "1111000101101100",
    "1110111110011001",
    "1110111000000011",
    "1110110011010011",
    "1110110000011110",
    "1110101111011110",
    "1110101111111011",
    "1110110001011001",
    "1110110011001101",
    "1110110100111001",
    "1110110110001101",
    "1110110111000001",
    "1110110111011011",
    "1110110111101100",
    "1110111000000100",
    "1110111000110101",
    "1110111010001001",
    "1110111011111111",
    "1110111110001101",
    "1111000000100111",
    "1111000010110100",
    "1111000100100100",
    "1111000101100101",
    "1111000101110001",
    "1111000101000101",
    "1111000011101010",
    "1111000001110001",
    "1110111111110011",
    "1110111110111101",
    "1111000001101011",
    "1111001010100110",
    "1111011011011110",
    "1111110011110110",
    "1111101111000101",
    "1111010001111000",
    "1110111001010011",
    "1110101001000100",
    "1110100010001111",
    "1110100011001111",
    "1110101000110010",
    "1110101111010010",
    "1110110100001000",
    "1110110110001101",
    "1110110101101010",
    "1110110011011100",
    "1110110000101011",
    "1110101101111101",
    "1110101011011110",
    "1110101001000100",
    "1110100110100100",
    "1110100100000011",
    "1110100001111000",
    "1110100000010001",
    "1110011111010010",
    "1110011110101000",
    "1110011101111111",
    "1110011101010110",
    "1110011100111010",
    "1110011100111111",
    "1110011110000000",
    "1110100000010101",
    "1110100100010000",
    "1110101001111100",
    "1110110001100111",
    "1110111011011110",
    "1111000111010110",
    "1111010100011111",
    "1111100001011100",
    "1111101100010111",
    "1111110011101100",
    "1111110110100110",
    "1111110101011101",
    "1111110001110101",
    "1111101101111110",
    "1111101011111111",
    "1111101101000110",
    "1111110001001001",
    "1111110110111000",
    "1111111100011111",
    "1111111111101101",
    "1111111110111001",
    "1111111110110000",
    "1111111001110010",
    "1111110011001010",
    "1111101100000111",
    "1111100101110001",
    "1111100000111101",
    "1111011110010110",
    "1111011110010100",
    "1111100001000010",
    "1111100110001101",
    "1111101101001101",
    "1111110101000100",
    "1111111100110011",
    "1111111100010111",
    "1111110111000110",
    "1111110011100100",
    "1111110001100010",
    "1111110000100001",
    "1111101111110001",
    "1111101110100001",
    "1111101100001010",
    "1111101000001110",
    "1111100010100111",
    "1111011011100001",
    "1111010011010011",
    "1111001010100101",
    "1111000010000000",
    "1110111010011110",
    "1110110100110110",
    "1110110001111110",
    "1110110010010111",
    "1110110101111011",
    "1110111100000010",
    "1111000011100010",
    "1111001010111010",
    "1111010000101100",
    "1111010011111000",
    "1111010011111110",
    "1111010001001000",
    "1111001011111101",
    "1111000101001011",
    "1110111101100100",
    "1110110101111100",
    "1110101110111111",
    "1110101001010110",
    "1110100101100100",
    "1110100011111001",
    "1110100100011000",
    "1110100110110001",
    "1110101010100010",
    "1110101111000100",
    "1110110011101110",
    "1110110111110010",
    "1110111010100110",
    "1110111011100101",
    "1110111010010011",
    "1110110110101111",
    "1110110001010100",
    "1110101010111010",
    "1110100100100101",
    "1110011111100001",
    "1110011100101010",
    "1110011100100011",
    "1110011111010111",
    "1110100100111001",
    "1110101100101101",
    "1110110110010011",
    "1111000001000010",
    "1111001100001100",
    "1111010110111110",
    "1111100000011111",
    "1111100111111100",
    "1111101100101001",
    "1111101110010100",
    "1111101101000110",
    "1111101001011111",
    "1111100100011101",
    "1111011111000101",
    "1111011010100000",
    "1111010111100101",
    "1111010110110111",
    "1111011000100011",
    "1111011100010011",
    "1111100001011111",
    "1111100111010010",
    "1111101100101010",
    "1111110000100110",
    "1111110010001010",
    "1111110000101111",
    "1111101100000111",
    "1111100100101100",
    "1111011011010011",
    "1111010001000111",
    "1111000111010110",
    "1110111111001010",
    "1110111001010001",
    "1110110110000001",
    "1110110101011000",
    "1110110111001011",
    "1110111011000111",
    "1111000000111101",
    "1111001000100000",
    "1111010001010101",
    "1111011010111101",
    "1111100100100101",
    "1111101101011100",
    "1111110100110100",
    "1111111010001111",
    "1111111101101000",
    "1111111111000101",
    "1111111110111010",
    "1111111101011101",
    "1111111011000010",
    "1111110111111111",
    "1111110100100100",
    "1111110001000111",
    "1111101101110111",
    "1111101011000111",
    "1111101001000110",
    "1111101000000011",
    "1111101000001011",
    "1111101001100101",
    "1111101100001100",
    "1111101111110011",
    "1111110100000011",
    "1111111000100010",
    "1111111100110110",
    "1111111111001101",
    "1111111011111110",
    "1111111001100010",
    "1111111000000001",
    "1111110111100100",
    "1111111000010001",
    "1111111010000101",
    "1111111100110110",
    "1111111111101000",
    "1111111011110010",
    "1111110111110001",
    "1111110011110000",
    "1111101111111101",
    "1111101100101101",
    "1111101010100011",
    "1111101010000110",
    "1111101011111000",
    "1111110000000111",
    "1111110110100110",
    "1111111110101101",
    "1111111000010101",
    "1111101111011001",
    "1111100111000001",
    "1111011111010110",
    "1111011000010000",
    "1111010001100001",
    "1111001011000010",
    "1111000101001000",
    "1111000000001111",
    "1110111101000101",
    "1110111100010011",
    "1110111110001010",
    "1111000010100100",
    "1111001001000010",
    "1111010000110101",
    "1111011001000010",
    "1111100000111101",
    "1111100111111101",
    "1111101101110001",
    "1111110010010110",
    "1111110101110101",
    "1111111000011110",
    "1111111010100011",
    "1111111100010100",
    "1111111101111010",
    "1111111111011011",
    "1111111111001000",
    "1111111101111100",
    "1111111101001010",
    "1111111100111011",
    "1111111101010001",
    "1111111110000101",
    "1111111111000110",
    "1111111111111101",
    "1111111111100101",
    "1111111111111101",
    "1111111110110010",
    "1111111100111001",
    "1111111010100111",
    "1111111000011111",
    "1111110111000010",
    "1111110110110001",
    "1111111000000101",
    "1111111011010000",
    "1111111111100010",
    "1111111000011010",
    "1111101111011010",
    "1111100100101001",
    "1111011000001100",
    "1111001010011011",
    "1110111100000001",
    "1110101101111101",
    "1110100001011110",
    "1110010111100101",
    "1110010000111001",
    "1110001101011110",
    "1110001100110000",
    "1110001101110101",
    "1110001111111011",
    "1110010010100010",
    "1110010101100101",
    "1110011001010000",
    "1110011101101101",
    "1110100011000001",
    "1110101001000010",
    "1110101111011110",
    "1110110110000110",
    "1110111100110011",
    "1111000011100110",
    "1111001010100000",
    "1111010001011010",
    "1111011000000011",
    "1111011101110010",
    "1111100010001000",
    "1111100100101111",
    "1111100101101100",
    "1111100101010000",
    "1111100011110100",
    "1111100001110001",
    "1111011111001111",
    "1111011100001001",
    "1111011000001011",
    "1111010010111101",
    "1111001100011001",
    "1111000100101001",
    "1110111100010001",
    "1110110100000110",
    "1110101101000101",
    "1110101000000110",
    "1110100101101100",
    "1110100110001000",
    "1110101001010110",
    "1110101111000101",
    "1110110110111111",
    "1111000000101011",
    "1111001011101011",
    "1111010111011101",
    "1111100011010111",
    "1111101110101001",
    "1111111000101100",
    "1111111111000010",
    "1111111000110101",
    "1111110100101011",
    "1111110010010100",
    "1111110001010110",
    "1111110001011000",
    "1111110010000011",
    "1111110011001001",
    "1111110100100011",
    "1111110110010010",
    "1111111000100001",
    "1111111011100011",
    "1111111111101101",
    "1111111010101011",
    "1111110011101000",
    "1111101011011001",
    "1111100010100100",
    "1111011010000001",
    "1111010010100010",
    "1111001100110010",
    "1111001000111100",
    "1111000110110010",
    "1111000101111001",
    "1111000101110001",
    "1111000110001011",
    "1111000111000110",
    "1111001000110100",
    "1111001011101010",
    "1111001111111000",
    "1111010101100000",
    "1111011100010100",
    "1111100100000001",
    "1111101100010011",
    "1111110100111110",
    "1111111110000000",
    "1111111000100110",
    "1111101110111110",
    "1111100101010111",
    "1111011100001110",
    "1111010100001010",
    "1111001101101101",
    "1111001001000111",
    "1111000110011101",
    "1111000101011000",
    "1111000101011101",
    "1111000110001110",
    "1111000111010001",
    "1111001000011010",
    "1111001001011000",
    "1111001010000110",
    "1111001010010110",
    "1111001001110111",
    "1111001000011011",
    "1111000101111001",
    "1111000010010010",
    "1110111101111011",
    "1110111001010001",
    "1110110100111110",
    "1110110001101110",
    "1110110000000000",
    "1110110000000000",
    "1110110001011010",
    "1110110011101001",
    "1110110101111011",
    "1110110111100011",
    "1110111000000011",
    "1110110111010001",
    "1110110101011101",
    "1110110010111101",
    "1110110000001010",
    "1110101101011011",
    "1110101010110111",
    "1110101000100101",
    "1110100110100010",
    "1110100100101111",
    "1110100011010000",
    "1110100010010000",
    "1110100001111101",
    "1110100010101001",
    "1110100100100100",
    "1110101000010011",
    "1110101111011111",
    "1110111100001100",
    "1111001111110011",
    "1111101010000100",
    "1111110111010001",
    "1111011000001100",
    "1110111100111111",
    "1110101001000100",
    "1110011101111101",
    "1110011010101101",
    "1110011100110010",
    "1110100001001101",
    "1110100101100010",
    "1110101000101000",
    "1110101010010011",
    "1110101010111111",
    "1110101011011001",
    "1110101011111101",
    "1110101100100110",
    "1110101101010001",
    "1110101101110000",
    "1110101110000111",
    "1110101110101011",
    "1110101111101011",
    "1110110001000101",
    "1110110010100111",
    "1110110011111110",
    "1110110101000001",
    "1110110101111001",
    "1110110110110010",
    "1110110111111100",
    "1110111001101000",
    "1110111100010001",
    "1111000000101001",
    "1111000111101111",
    "1111010010000101",
    "1111011111011110",
    "1111101110011110",
    "1111111100101010",
    "1111111000101100",
    "1111110011111111",
    "1111110110001001",
    "1111111110011000",
    "1111110101011100",
    "1111101000010111",
    "1111011101001010",
    "1111010101110001",
    "1111010010110001",
    "1111010011110110",
    "1111010111111001",
    "1111011101110000",
    "1111100100011100",
    "1111101011001000",
    "1111110001000001",
    "1111110101010111",
    "1111110111011111",
    "1111110111000111",
    "1111110100101000",
    "1111110000111111",
    "1111101101100111",
    "1111101100000010",
    "1111101101011000",
    "1111110010000010",
    "1111111001101100",
    "1111111100100000",
    "1111110001110010",
    "1111100111001110",
    "1111011101110000",
    "1111010110000110",
    "1111010000110011",
    "1111001110010010",
    "1111001110110000",
    "1111010010001010",
    "1111010111111100",
    "1111011111001111",
    "1111100110111000",
    "1111101101110001",
    "1111110011001110",
    "1111110111000011",
    "1111111001011111",
    "1111111010111100",
    "1111111011101001",
    "1111111011100101",
    "1111111010010100",
    "1111110111001110",
    "1111110001110100",
    "1111101001111001",
    "1111011111110000",
    "1111010100001011",
    "1111001000010011",
    "1110111101010001",
    "1110110100000000",
    "1110101100111000",
    "1110100111110100",
    "1110100100001010",
    "1110100000111001",
    "1110011101000100",
    "1110010111110100",
    "1110010000110101",
    "1110001000010000",
    "1101111110101110",
    "1101110101001101",
    "1101101100101110",
    "1101100110010010",
    "1101100010011101",
    "1101100001101011",
    "1101100100000001",
    "1101101001011101",
    "1101110001111000",
    "1101111100111111",
    "1110001010001100",
    "1110011000110100",
    "1110100111110010",
    "1110110110001001",
    "1111000011000101",
    "1111001110001111",
    "1111010111110100",
    "1111100000100001",
    "1111101001001000",
    "1111110010010001",
    "1111111100001111",
    "1111111001001000",
    "1111101110011001",
    "1111100100001010",
    "1111011010110111",
    "1111010010111001",
    "1111001100010100",
    "1111000111001101",
    "1111000011101010",
    "1111000001111000",
    "1111000010000000",
    "1111000100010010",
    "1111001000110100",
    "1111001111101110",
    "1111011001000010",
    "1111100100011111",
    "1111110001100100",
    "1111111111011100",
    "1111110010111110",
    "1111100110111110",
    "1111011101101101",
    "1111010111111100",
    "1111010101110111",
    "1111010111000011",
    "1111011010101010",
    "1111011111101100",
    "1111100101010011",
    "1111101010111001",
    "1111110000010010",
    "1111110101011000",
    "1111111010000110",
    "1111111110001100",
    "1111111110101110",
    "1111111101000100",
    "1111111100111110",
    "1111111110010101",
    "1111111111001011",
    "1111111100001010",
    "1111111000111111",
    "1111110101111000",
    "1111110010110110",
    "1111101111110100",
    "1111101100101100",
    "1111101001101000",
    "1111100110111001",
    "1111100100110110",
    "1111100011110100",
    "1111100100000001",
    "1111100101011010",
    "1111100111110001",
    "1111101010101011",
    "1111101101110000",
    "1111110000101100",
    "1111110011010100",
    "1111110101100111",
    "1111110111100101",
    "1111111001001110",
    "1111111010010111",
    "1111111010110000",
    "1111111010001101",
    "1111111000101110",
    "1111110110101000",
    "1111110100011111",
    "1111110010111100",
    "1111110010100000",
    "1111110011011001",
    "1111110101011110",
    "1111111000011001",
    "1111111011110000",
    "1111111111001010",
    "1111111101011111",
    "1111111010010101",
    "1111110111001111",
    "1111110100001101",
    "1111110001001010",
    "1111101110001011",
    "1111101011011010",
    "1111101001000001",
    "1111100111001110",
    "1111100110001101",
    "1111100110000110",
    "1111100110111111",
    "1111101000110011",
    "1111101011011011",
    "1111101110101001",
    "1111110010001101",
    "1111110101110011",
    "1111111001001001",
    "1111111011111110",
    "1111111110001000",
    "1111111111100011",
    "1111111111101001",
    "1111111111011011",
    "1111111111101010",
    "1111111111100101",
    "1111111110010001",
    "1111111100001100",
    "1111111001001010",
    "1111110101001000",
    "1111110000001111",
    "1111101010110000",
    "1111100101001000",
    "1111011111111000",
    "1111011011100101",
    "1111011000110101",
    "1111011000000011",
    "1111011001100010",
    "1111011101010010",
    "1111100010111110",
    "1111101010000001",
    "1111110001101010",
    "1111111001001000",
    "1111111111101110",
    "1111111010111101",
    "1111110111001100",
    "1111110100111010",
    "1111110011111011",
    "1111110011111100",
    "1111110100101110",
    "1111110110000001",
    "1111110111101010",
    "1111111001011110",
    "1111111011010100",
    "1111111101000011",
    "1111111110100011",
    "1111111111110011",
    "1111111111000110",
    "1111111110000011",
    "1111111100101100",
    "1111111010110011",
    "1111111000001010",
    "1111110100110101",
    "1111110000111110",
    "1111101100111001",
    "1111101000111110",
    "1111100101011101",
    "1111100010100010",
    "1111100000001101",
    "1111011110010110",
    "1111011100110111",
    "1111011011110010",
    "1111011011010001",
    "1111011011100101",
    "1111011101000010",
    "1111011111101100",
    "1111100011011111",
    "1111100111111111",
    "1111101100101010",
    "1111110000111010",
    "1111110100001010",
    "1111110101111110",
    "1111110110000111",
    "1111110100100000",
    "1111110001001011",
    "1111101100010010",
    "1111100110000110",
    "1111011110111101",
    "1111010111010000",
    "1111001111010100",
    "1111000111100011",
    "1111000000010100",
    "1110111001111001",
    "1110110100100010",
    "1110110000011100",
    "1110101101110000",
    "1110101100011011",
    "1110101100011011",
    "1110101101101011",
    "1110110000001000",
    "1110110011110110",
    "1110111000111001",
    "1110111111010110",
    "1111000111001001",
    "1111010000000011",
    "1111011001101000",
    "1111100011001011",
    "1111101011111110",
    "1111110011011000",
    "1111111000111011",
    "1111111100100000",
    "1111111110010001",
    "1111111110100111",
    "1111111110000001",
    "1111111100111001",
    "1111111011011101",
    "1111111001101110",
    "1111110111100001",
    "1111110100100111",
    "1111110000111000",
    "1111101100011101",
    "1111100111101010",
    "1111100011000001",
    "1111011111000000",
    "1111011011110011",
    "1111011001011011",
    "1111010111100101",
    "1111010101110111",
    "1111010011111110",
    "1111010001110001",
    "1111001111011001",
    "1111001101000101",
    "1111001011001110",
    "1111001010000001",
    "1111001001100011",
    "1111001001110100",
    "1111001010100101",
    "1111001011101011",
    "1111001100111101",
    "1111001110010001",
    "1111001111101000",
    "1111010001000011",
    "1111010010101011",
    "1111010100100100",
    "1111010110110110",
    "1111011001101101",
    "1111011101010010",
    "1111100001110100",
    "1111100111100101",
    "1111101110110010",
    "1111110111011110",
    "1111111110100001",
    "1111110011101110",
    "1111101000110011",
    "1111011110100001",
    "1111010101011011",
    "1111001101110111",
    "1111000111101100",
    "1111000010100111",
    "1110111110010100",
    "1110111010100110",
    "1110110111100111",
    "1110110101100010",
    "1110110100101010",
    "1110110100111110",
    "1110110110001101",
    "1110110111110101",
    "1110111001010011",
    "1110111010001001",
    "1110111010001111",
    "1110111001101111",
    "1110111000110101",
    "1110110111111001",
    "1110110110111110",
    "1110110110001001",
    "1110110101010111",
    "1110110100100000",
    "1110110011100110",
    "1110110010101011",
    "1110110001111000",
    "1110110001010101",
    "1110110001001111",
    "1110110001100100",
    "1110110010011100",
    "1110110011111000",
    "1110110110100100",
    "1110111100010111",
    "1111000111110100",
    "1111011010100000",
    "1111110100001000",
    "1111101110000101",
    "1111010000101110",
    "1110111000100010",
    "1110101001001100",
    "1110100011101010",
    "1110100110000001",
    "1110101100101011",
    "1110110011101100",
    "1110111000011010",
    "1110111001111001",
    "1110111000101000",
    "1110110101111110",
    "1110110011010011",
    "1110110001010101",
    "1110110000001010",
    "1110101111010110",
    "1110101110010111",
    "1110101101000000",
    "1110101011011011",
    "1110101001111001",
    "1110101000100000",
    "1110100111001110",
    "1110100110000000",
    "1110100101000000",
    "1110100100100111",
    "1110100101001110",
    "1110100111001011",
    "1110101010100110",
    "1110101111011010",
    "1110110101100000",
    "1110111100101000",
    "1111000100011111",
    "1111001100110010",
    "1111010101000000",
    "1111011100100101",
    "1111100011000011",
    "1111101000001000",
    "1111101011111010",
    "1111101110110111",
    "1111110001101001",
    "1111110100110111",
    "1111111000110100",
    "1111111101001100",
    "1111111110110111",
    "1111111100100110",
    "1111111100111001",
    "1111111111111011",
    "1111111010011000",
    "1111110011011110",
    "1111101100011110",
    "1111100110011101",
    "1111100010000110",
    "1111011111110011",
    "1111011111100100",
    "1111100001010101",
    "1111100101000101",
    "1111101010110011",
    "1111110010010111",
    "1111111011010011",
    "1111111011010011",
    "1111110010101101",
    "1111101100000010",
    "1111101000000010",
    "1111100110110111",
    "1111100111111000",
    "1111101001111100",
    "1111101011100111",
    "1111101011110010",
    "1111101001110100",
    "1111100101101010",
    "1111011111101011",
    "1111011000100010",
    "1111010000110110",
    "1111001001010001",
    "1111000010010101",
    "1110111100100001",
    "1110111000011110",
    "1110110110110001",
    "1110110111101101",
    "1110111011011001",
    "1111000001010000",
    "1111001000010101",
    "1111001111001101",
    "1111010100100111",
    "1111010111011111",
    "1111010111011011",
    "1111010100100100",
    "1111001111011111",
    "1111001000111100",
    "1111000001100010",
    "1110111001101111",
    "1110110001101110",
    "1110101001110111",
    "1110100010100100",
    "1110011100011011",
    "1110011000001001",
    "1110010110010000",
    "1110010110111110",
    "1110011010000100",
    "1110011110111111",
    "1110100100110111",
    "1110101010111100",
    "1110110000011111",
    "1110110101000001",
    "1110111000010001",
    "1110111010000110",
    "1110111010011001",
    "1110111001001100",
    "1110110110101000",
    "1110110011000011",
    "1110101111000010",
    "1110101011011011",
    "1110101001000110",
    "1110101000111100",
    "1110101011100011",
    "1110110001000101",
    "1110111001010001",
    "1111000011010010",
    "1111001110000111",
    "1111011000101000",
    "1111100001111000",
    "1111101001010011",
    "1111101110100111",
    "1111110001110101",
    "1111110011000100",
    "1111110010011110",
    "1111110000001011",
    "1111101100011110",
    "1111100111101110",
    "1111100010100001",
    "1111011101010110",
    "1111011000110000",
    "1111010101000110",
    "1111010010011100",
    "1111010000101011",
    "1111001111100100",
    "1111001110111010",
    "1111001110100110",
    "1111001110100001",
    "1111001110101110",
    "1111001111001101",
    "1111001111111011",
    "1111010000110101",
    "1111010001111000",
    "1111010011000011",
    "1111010100011101",
    "1111010110001101",
    "1111011000010000",
    "1111011010100000",
    "1111011100101011",
    "1111011110011111",
    "1111011111110000",
    "1111100000011001",
    "1111100000101011",
    "1111100000111000",
    "1111100001010111",
    "1111100010010111",
    "1111100011111110",
    "1111100110001000",
    "1111101000101101",
    "1111101011100010",
    "1111101110011111",
    "1111110001011011",
    "1111110100001000",
    "1111110110011110",
    "1111111000010010",
    "1111111001100110",
    "1111111010100001",
    "1111111011010011",
    "1111111100010001",
    "1111111101100111",
    "1111111111010000",
    "1111111110111101",
    "1111111101100100",
    "1111111100111110",
    "1111111101100000",
    "1111111111001100",
    "1111111110001011",
    "1111111011001001",
    "1111111000001011",
    "1111110101101010",
    "1111110011101111",
    "1111110010011001",
    "1111110001011100",
    "1111110000110010",
    "1111110000011011",
    "1111110000011110",
    "1111110001000101",
    "1111110010011111",
    "1111110100110011",
    "1111111000000111",
    "1111111100011110",
    "1111111110001001",
    "1111110111111000",
    "1111110000111010",
    "1111101001100110",
    "1111100010010111",
    "1111011011110011",
    "1111010110011111",
    "1111010010110001",
    "1111010000111011",
    "1111010000111101",
    "1111010010100010",
    "1111010101010000",
    "1111011000100000",
    "1111011011101111",
    "1111011110011111",
    "1111100000011111",
    "1111100001100010",
    "1111100001101100",
    "1111100001000011",
    "1111011111110110",
    "1111011110010001",
    "1111011100101101",
    "1111011011100001",
    "1111011011001100",
    "1111011100000100",
    "1111011110011001",
    "1111100010001010",
    "1111100111000111",
    "1111101100110011",
    "1111110010101100",
    "1111111000010110",
    "1111111101011010",
    "1111111110010000",
    "1111111010110010",
    "1111111000001000",
    "1111110110010010",
    "1111110101010001",
    "1111110101000101",
    "1111110101101010",
    "1111110110111001",
    "1111111000100101",
    "1111111010100101",
    "1111111100110100",
    "1111111111010010",
    "1111111101110001",
    "1111111010001110",
    "1111110101110000",
    "1111110000001110",
    "1111101001100110",
    "1111100001111000",
    "1111011001000100",
    "1111001111001000",
    "1111000100001110",
    "1110111000101111",
    "1110101101010111",
    "1110100010111000",
    "1110011001111010",
    "1110010010111001",
    "1110001101111011",
    "1110001010111000",
    "1110001001100011",
    "1110001001110101",
    "1110001011111000",
    "1110010000000011",
    "1110010110100101",
    "1110011111100110",
    "1110101010110000",
    "1110110111010000",
    "1111000011111000",
    "1111001111010001",
    "1111011000001110",
    "1111011110000101",
    "1111100000110101",
    "1111100000111101",
    "1111011111010010",
    "1111011100101101",
    "1111011001110000",
    "1111010110110001",
    "1111010011110100",
    "1111010000110101",
    "1111001101101000",
    "1111001010000110",
    "1111000110000011",
    "1111000001011010",
    "1110111100001001",
    "1110110110010101",
    "1110110000011001",
    "1110101010110111",
    "1110100110011111",
    "1110100011110100",
    "1110100011010000",
    "1110100100111001",
    "1110101000101010",
    "1110101110010111",
    "1110110101111001",
    "1110111111001010",
    "1111001001110111",
    "1111010101100100",
    "1111100001011111",
    "1111101100101100",
    "1111110110010100",
    "1111111101101100",
    "1111111101010100",
    "1111111010011110",
    "1111111001000101",
    "1111111000011011",
    "1111110111111001",
    "1111110111010010",
    "1111110110110100",
    "1111110110111111",
    "1111111000011110",
    "1111111011111011",
    "1111111110001101",
    "1111110101111100",
    "1111101011101000",
    "1111100000001101",
    "1111010100111011",
    "1111001011001001",
    "1111000011111011",
    "1110111111110110",
    "1110111110110001",
    "1111000000000101",
    "1111000010110001",
    "1111000110000001",
    "1111001001001100",
    "1111001100001001",
    "1111001110111101",
    "1111010001111000",
    "1111010101000110",
    "1111011000101111",
    "1111011100101101",
    "1111100000111000",
    "1111100101001011",
    "1111101001101000",
    "1111101110011001",
    "1111110011101001",
    "1111111001100010",
    "1111111111111011",
    "1111111000111111",
    "1111110001111110",
    "1111101011010101",
    "1111100101100101",
    "1111100001001000",
    "1111011110001101",
    "1111011100110000",
    "1111011100011001",
    "1111011100100101",
    "1111011100100110",
    "1111011011110101",
    "1111011001111001",
    "1111010110101010",
    "1111010010010101",
    "1111001101011100",
    "1111001000100010",
    "1111000100001010",
    "1111000000011111",
    "1110111101100001",
    "1110111010111101",
    "1110111000100111",
    "1110110110010101",
    "1110110100010010",
    "1110110010101110",
    "1110110001110100",
    "1110110001100110",
    "1110110001110011",
    "1110110010000011",
    "1110110001111001",
    "1110110001000111",
    "1110101111100100",
    "1110101101011011",
    "1110101010110010",
    "1110100111110101",
    "1110100100101010",
    "1110100001010111",
    "1110011110000010",
    "1110011010111000",
    "1110011000001011",
    "1110010110010010",
    "1110010101100000",
    "1110010110000100",
    "1110011000001001",
    "1110011011101011",
    "1110100000101001",
    "1110100111010000",
    "1110110000010001",
    "1110111101000000",
    "1111001110101000",
    "1111100101011000",
    "1111111111110100",
    "1111100011100110",
    "1111001001010001",
    "1110110100001011",
    "1110100110011111",
    "1110100000011110",
    "1110100000101110",
    "1110100100110100",
    "1110101010001011",
    "1110101110110110",
    "1110110010000000",
    "1110110011100111",
    "1110110100010010",
    "1110110100101110",
    "1110110101010010",
    "1110110110001000",
    "1110110111001011",
    "1110111000001100",
    "1110111001001011",
    "1110111010000100",
    "1110111010110101",
    "1110111011011000",
    "1110111011100101",
    "1110111011011011",
    "1110111011000010",
    "1110111010101000",
    "1110111010100101",
    "1110111011011011",
    "1110111101111111",
    "1111000011011101",
    "1111001100101101",
    "1111011001101010",
    "1111101000111100",
    "1111111000000010",
    "1111111100000001",
    "1111110101111001",
    "1111110110111000",
    "1111111110011110",
    "1111110101011000",
    "1111100111101010",
    "1111011011001010",
    "1111010010000011",
    "1111001101001111",
    "1111001100101101",
    "1111001111101001",
    "1111010101000000",
    "1111011011101111",
    "1111100011000000",
    "1111101010000011",
    "1111110000000111",
    "1111110100100001",
    "1111110110110001",
    "1111110110111000",
    "1111110101011001",
    "1111110011011001",
    "1111110010000010",
    "1111110010010100",
    "1111110100110100",
    "1111111001100101",
    "1111111111101100",
    "1111110111101111",
    "1111101111010010",
    "1111100111000110",
    "1111011111111000",
    "1111011010001110",
    "1111010110100111",
    "1111010101010111",
    "1111010110011101",
    "1111011001101010",
    "1111011110011001",
    "1111100100000000",
    "1111101001110000",
    "1111101111001000",
    "1111110011111110",
    "1111111000010000",
    "1111111100000001",
    "1111111111001100",
    "1111111110011101",
    "1111111101011111",
    "1111111110100010",
    "1111111101110001",
    "1111110111000000",
    "1111101100111111",
    "1111100000000101",
    "1111010001001010",
    "1111000001100010",
    "1110110010101011",
    "1110100101110110",
    "1110011100000010",
    "1110010101100101",
    "1110010010001111",
    "1110010001000011",
    "1110010000110101",
    "1110010000010001",
    "1110001110010010",
    "1110001010010100",
    "1110000100010111",
    "1101111101000100",
    "1101110101011011",
    "1101101110101001",
    "1101101001100010",
    "1101100110100111",
    "1101100110000000",
    "1101100111100111",
    "1101101011010001",
    "1101110001000000",
    "1101111001000001",
    "1110000011101001",
    "1110010001000101",
    "1110100001001010",
    "1110110011001101",
    "1111000110001000",
    "1111011000101111",
    "1111101010000001",
    "1111111001001001",
    "1111111010001111",
    "1111110000001111",
    "1111101000100001",
    "1111100010101111",
    "1111011110100100",
    "1111011011101011",
    "1111011001110100",
    "1111011000110101",
    "1111011000101100",
    "1111011001011000",
    "1111011010111101",
    "1111011101100001",
    "1111100001000000",
    "1111100101010111",
    "1111101010010011",
    "1111101111011100",
    "1111110100010011",
    "1111111000011001",
    "1111111011011111",
    "1111111101100111",
    "1111111110111111",
    "1111111111111101",
    "1111111110111011",
    "1111111101100101",
    "1111111011110100",
    "1111111001101111",
    "1111110111100010",
    "1111110101011000",
    "1111110011011001",
    "1111110001100110",
    "1111101111111110",
    "1111101110100110",
    "1111101101100110",
    "1111101101001100",
    "1111101101011101",
    "1111101110011010",
    "1111101111110101",
    "1111110001011011",
    "1111110010110111",
    "1111110011111010",
    "1111110100011111",
    "1111110100100101",
    "1111110100010100",
    "1111110011110011",
    "1111110011001111",
    "1111110010110010",
    "1111110010100011",
    "1111110010100011",
    "1111110010110000",
    "1111110011000000",
    "1111110011001001",
    "1111110010111110",
    "1111110010010011",
    "1111110001000101",
    "1111101111001111",
    "1111101100110110",
    "1111101010000010",
    "1111100110111111",
    "1111100100000110",
    "1111100001110000",
    "1111100000011001",
    "1111100000010101",
    "1111100001111000",
    "1111100101000001",
    "1111101001101011",
    "1111101111101110",
    "1111110110111000",
    "1111111110110100",
    "1111111000110011",
    "1111110000100111",
    "1111101001001001",
    "1111100010111110",
    "1111011110100001",
    "1111011100000101",
    "1111011011110010",
    "1111011101101000",
    "1111100001011100",
    "1111100110111101",
    "1111101101101110",
    "1111110101000100",
    "1111111100001110",
    "1111111101100100",
    "1111111001000010",
    "1111110110100101",
    "1111110110010100",
    "1111111000000101",
    "1111111011011001",
    "1111111111110000",
    "1111111011011100",
    "1111110110110010",
    "1111110010101100",
    "1111101111011101",
    "1111101101001111",
    "1111101100000011",
    "1111101011110010",
    "1111101100010011",
    "1111101101010011",
    "1111101110100010",
    "1111101111101111",
    "1111110000101011",
    "1111110001001000",
    "1111110000111101",
    "1111110000001000",
    "1111101110101110",
    "1111101100111010",
    "1111101011000001",
    "1111101001011111",
    "1111101000101111",
    "1111101001001010",
    "1111101010111101",
    "1111101110001000",
    "1111110010100001",
    "1111110111101101",
    "1111111101001110",
    "1111111101011101",
    "1111111000110011",
    "1111110101000111",
    "1111110010100011",
    "1111110001001001",
    "1111110000111011",
    "1111110001110110",
    "1111110011111010",
    "1111110111000001",
    "1111111011000010",
    "1111111111101011",
    "1111111011011010",
    "1111110110110010",
    "1111110010111100",
    "1111110000001011",
    "1111101110100111",
    "1111101110000101",
    "1111101110001111",
    "1111101110101001",
    "1111101110111100",
    "1111101110111011",
    "1111101110100000",
    "1111101101110011",
    "1111101100111110",
    "1111101100001011",
    "1111101011100001",
    "1111101011000111",
    "1111101010111100",
    "1111101011000000",
    "1111101011001110",
    "1111101011100010",
    "1111101011110100",
    "1111101011111110",
    "1111101011111000",
    "1111101011011000",
    "1111101010010110",
    "1111101000100101",
    "1111100101111110",
    "1111100010011001",
    "1111011101111010",
    "1111011000101000",
    "1111010010110001",
    "1111001100100000",
    "1111000110001001",
    "1111000000000010",
    "1110111010100011",
    "1110110101111001",
    "1110110010001011",
    "1110101111011001",
    "1110101101010110",
    "1110101011110111",
    "1110101010111100",
    "1110101010111010",
    "1110101100010111",
    "1110110000000101",
    "1110110110100101",
    "1111000000000000",
    "1111001011110000",
    "1111011000101000",
    "1111100100111100",
    "1111101111001011",
    "1111110110001001",
    "1111111001100011",
    "1111111001110110",
    "1111111000000001",
    "1111110101001001",
    "1111110010000101",
    "1111101111001101",
    "1111101100100001",
    "1111101001101110",
    "1111100110100000",
    "1111100010101111",
    "1111011110101000",
    "1111011010101010",
    "1111010111011010",
    "1111010101010011",
    "1111010100100100",
    "1111010100111100",
    "1111010110000011",
    "1111010111010011",
    "1111011000010000",
    "1111011000100111",
    "1111011000010001",
    "1111010111011010",
    "1111010110001001",
    "1111010100110100",
    "1111010011101001",
    "1111010010111011",
    "1111010010110001",
    "1111010011001010",
    "1111010011111000",
    "1111010100100010",
    "1111010100100101",
    "1111010011100001",
    "1111010001000000",
    "1111001101000000",
    "1111001000000100",
    "1111000010111001",
    "1110111110100110",
    "1110111100000100",
    "1110111100000010",
    "1110111110110110",
    "1111000100101001",
    "1111001101010001",
    "1111011000011010",
    "1111100101100000",
    "1111110011110110",
    "1111111101101100",
    "1111110000011000",
    "1111100101001110",
    "1111011100111000",
    "1111010111011000",
    "1111010100000001",
    "1111010001110000",
    "1111001111010110",
    "1111001100000001",
    "1111000111100111",
    "1111000010100110",
    "1110111101111011",
    "1110111010100000",
    "1110111000101101",
    "1110111000011101",
    "1110111001000110",
    "1110111001101101",
    "1110111001100011",
    "1110111000010000",
    "1110110101110110",
    "1110110010101001",
    "1110101111001000",
    "1110101011110000",
    "1110101000110101",
    "1110100110101000",
    "1110100101010011",
    "1110100100111100",
    "1110100101100101",
    "1110100111001000",
    "1110101001010110",
    "1110101100000010",
    "1110101110111000",
    "1110110001100110",
    "1110110100000110",
    "1110110111001101",
    "1110111101000000",
    "1111001000010001",
    "1111011010110010",
    "1111110100010000",
    "1111101110001010",
    "1111010001000101",
    "1110111001010000",
    "1110101010001110",
    "1110100100110110",
    "1110100111001001",
    "1110101101101001",
    "1110110100101001",
    "1110111001101011",
    "1110111100000100",
    "1110111100001010",
    "1110111011000110",
    "1110111001110111",
    "1110111000110000",
    "1110110111101000",
    "1110110110000100",
    "1110110011110001",
    "1110110000111000",
    "1110101101111111",
    "1110101011101000",
    "1110101010000110",
    "1110101001010000",
    "1110101000111001",
    "1110101000111010",
    "1110101001011000",
    "1110101010011110",
    "1110101100010110",
    "1110101111001100",
    "1110110011000101",
    "1110111000001011",
    "1110111110011111",
    "1111000101110110",
    "1111001101110000",
    "1111010101100111",
    "1111011100101010",
    "1111100010010111",
    "1111100110011101",
    "1111101001001011",
    "1111101011001000",
    "1111101101000110",
    "1111101111101111",
    "1111110011010101",
    "1111110111100101",
    "1111111011101010",
    "1111111110100001",
    "1111111111010001",
    "1111111101101001",
    "1111111001111100",
    "1111110100111110",
    "1111101111101001",
    "1111101010110010",
    "1111100111000010",
    "1111100100110011",
    "1111100100010101",
    "1111100101110001",
    "1111101001000110",
    "1111101110010110",
    "1111110101010100",
    "1111111101100011",
    "1111111001100011",
    "1111110000110110",
    "1111101000111111",
    "1111100010100100",
    "1111011110000000",
    "1111011011011001",
    "1111011010100010",
    "1111011010111010",
    "1111011011111000",
    "1111011100110010",
    "1111011101000100",
    "1111011100100011",
    "1111011011010100",
    "1111011001101010",
    "1111010111111110",
    "1111010110011000",
    "1111010100111001",
    "1111010011010101",
    "1111010001011110",
    "1111001111001101",
    "1111001100101000",
    "1111001001110111",
    "1111000111000110",
    "1111000100100010",
    "1111000010001101",
    "1111000000001000",
    "1110111110010001",
    "1110111100100001",
    "1110111010111100",
    "1110111001011011",
    "1110110111111111",
    "1110110110100010",
    "1110110100110110",
    "1110110010110001",
    "1110110000001000",
    "1110101100110111",
    "1110101001000110",
    "1110100101001000",
    "1110100001011010",
    "1110011110011100",
    "1110011100100011",
    "1110011011110010",
    "1110011100000001",
    "1110011100111111",
    "1110011110011110",
    "1110100000011100",
    "1110100011000000",
    "1110100110010101",
    "1110101010100000",
    "1110101111011111",
    "1110110101000000",
    "1110111010101010",
    "1111000000000011",
    "1111000100111100",
    "1111001001000110",
    "1111001100010111",
    "1111001110110101",
    "1111010000011100",
    "1111010001010100",
    "1111010001100001",
    "1111010001001111",
    "1111010000100100",
    "1111001111110000",
    "1111001110111111",
    "1111001110100001",
    "1111001110100011",
    "1111001111010001",
    "1111010000101001",
    "1111010010101111",
    "1111010101011010",
    "1111011000011101",
    "1111011011100101",
    "1111011110011100",
    "1111100000110001",
    "1111100010001101",
    "1111100010100100",
    "1111100001110001",
    "1111011111111011",
    "1111011101001100",
    "1111011001110111",
    "1111010110010101",
    "1111010010111001",
    "1111001111111000",
    "1111001101011110",
    "1111001011110101",
    "1111001011000010",
    "1111001011001001",
    "1111001100001001",
    "1111001101111010",
    "1111010000001111",
    "1111010010111101",
    "1111010101101111",
    "1111011000011010",
    "1111011010110100",
    "1111011101000000",
    "1111011111000111",
    "1111100001010010",
    "1111100011101111",
    "1111100110101000",
    "1111101001111100",
    "1111101101101001",
    "1111110001101001",
    "1111110101110011",
    "1111111001110011",
    "1111111101010100",
    "1111111111111000",
    "1111111110111101",
    "1111111111100100",
    "1111111110000101",
    "1111111010011100",
    "1111110110010000",
    "1111110010010010",
    "1111101111001101",
    "1111101101001111",
    "1111101100010011",
    "1111101100001011",
    "1111101100101010",
    "1111101101101101",
    "1111101111011011",
    "1111110001111110",
    "1111110101010101",
    "1111111001010001",
    "1111111101010111",
    "1111111110111011",
    "1111111100001011",
    "1111111010101110",
    "1111111010110010",
    "1111111100010000",
    "1111111110110110",
    "1111111101111011",
    "1111111010110100",
    "1111111000011010",
    "1111110111010001",
    "1111110111101110",
    "1111111001111010",
    "1111111101101101",
    "1111111101000101",
    "1111110110110101",
    "1111101111111001",
    "1111101000100111",
    "1111100001011001",
    "1111011010101010",
    "1111010100110100",
    "1111010000001111",
    "1111001101001100",
    "1111001011101111",
    "1111001011110010",
    "1111001101000101",
    "1111001111001101",
    "1111010001110000",
    "1111010100001110",
    "1111010110010011",
    "1111010111110001",
    "1111011000100010",
    "1111011000101100",
    "1111011000100011",
    "1111011000100011",
    "1111011001001100",
    "1111011010110101",
    "1111011101110011",
    "1111100010000110",
    "1111100111100000",
    "1111101101100100",
    "1111110011101111",
    "1111111001100010",
    "1111111110101010",
    "1111111101000001",
    "1111111001100110",
    "1111110110111011",
    "1111110101000000",
    "1111110011110011",
    "1111110011010100",
    "1111110011100001",
    "1111110100010101",
    "1111110101100101",
    "1111110111001110",
    "1111111001010111",
    "1111111100010110",
    "1111111111010010",
    "1111111001000101",
    "1111110000101101",
    "1111100110001011",
    "1111011001111010",
    "1111001100101011",
    "1110111111010110",
    "1110110010111101",
    "1110101000011110",
    "1110100000100100",
    "1110011011011101",
    "1110011001000001",
    "1110011000110100",
    "1110011010001100",
    "1110011100100110",
    "1110011111101011",
    "1110100011010011",
    "1110100111100010",
    "1110101100011001",
    "1110110001110110",
    "1110110111110010",
    "1110111101111101",
    "1111000100000001",
    "1111001001101010",
    "1111001110101011",
    "1111010010111110",
    "1111010110100000",
    "1111011001000111",
    "1111011010100110",
    "1111011010101000",
    "1111011000111010",
    "1111010101011111",
    "1111010000011010",
    "1111001001110000",
    "1111000001110000",
    "1110111000101101",
    "1110101111001111",
    "1110100110001110",
    "1110011110100110",
    "1110011001001011",
    "1110010110010110",
    "1110010110001101",
    "1110011000011011",
    "1110011100101011",
    "1110100010101111",
    "1110101010101010",
    "1110110100010101",
    "1110111111011001",
    "1111001011000111",
    "1111010110100111",
    "1111100001000011",
    "1111101001110100",
    "1111110000101000",
    "1111110101100100",
    "1111111000111001",
    "1111111011000000",
    "1111111100001101",
    "1111111100110000",
    "1111111100110101",
    "1111111100110001",
    "1111111100101100",
    "1111111100100110",
    "1111111100000010",
    "1111111010011011",
    "1111110111000110",
    "1111110001101001",
    "1111101010000110",
    "1111100001000011",
    "1111010111100101",
    "1111001110110110",
    "1111000111111111",
    "1111000011101100",
    "1111000001111110",
    "1111000010011010",
    "1111000100000001",
    "1111000101110010",
    "1111000110111001",
    "1111000110111110",
    "1111000110001110",
    "1111000101010000",
    "1111000100101100",
    "1111000100110111",
    "1111000101111011",
    "1111000111110001",
    "1111001010010110",
    "1111001101110011",
    "1111010010011100",
    "1111011000100010",
    "1111100000001010",
    "1111101001000000",
    "1111110010010111",
    "1111111011010111",
    "1111111100101011",
    "1111110110001001",
    "1111110000110011",
    "1111101100001001",
    "1111100111100000",
    "1111100010011100",
    "1111011100111100",
    "1111010111010011",
    "1111010010000110",
    "1111001101110111",
    "1111001010110111",
    "1111001001000110",
    "1111001000010000",
    "1111000111111100",
    "1111000111110010",
    "1111000111010110",
    "1111000110011010",
    "1111000100110110",
    "1111000010101001",
    "1110111111111101",
    "1110111100111101",
    "1110111001110111",
    "1110110110111001",
    "1110110100010011",
    "1110110010010000",
    "1110110000110001",
    "1110101111110101",
    "1110101111001100",
    "1110101110100100",
    "1110101101101011",
    "1110101100001110",
    "1110101010000100",
    "1110100111001110",
    "1110100011110110",
    "1110100000001111",
    "1110011100110011",
    "1110011001111111",
    "1110011000001000",
    "1110010111011011",
    "1110010111110111",
    "1110011001010101",
    "1110011011100101",
    "1110011110010100",
    "1110100001011100",
    "1110100100110011",
    "1110101000011101",
    "1110101100100110",
    "1110110010000101",
    "1110111010011011",
    "1111000111011000",
    "1111011010000110",
    "1111110010010111",
    "1111110001100111",
    "1111010101001101",
    "1110111100001100",
    "1110101001110111",
    "1110011111110000",
    "1110011101011001",
    "1110100000110110",
    "1110100111010011",
    "1110101110001111",
    "1110110100000000",
    "1110110111110101",
    "1110111001111101",
    "1110111010111000",
    "1110111011001001",
    "1110111011000010",
    "1110111010110100",
    "1110111010011110",
    "1110111010001111",
    "1110111010010001",
    "1110111010101101",
    "1110111011100000",
    "1110111100010111",
    "1110111101001001",
    "1110111101100110",
    "1110111101110011",
    "1110111101111010",
    "1110111110010001",
    "1110111111010010",
    "1111000001110000",
    "1111000110011011",
    "1111001101111010",
    "1111011000001011",
    "1111100100010010",
    "1111110000011111",
    "1111111010011110",
    "1111111111111010",
    "1111111111111000",
    "1111111001111000",
    "1111101111010100",
    "1111100010010101",
    "1111010101011101",
    "1111001010110010",
    "1111000011101100",
    "1111000000101001",
    "1111000001010111",
    "1111000101001000",
    "1111001011001010",
    "1111010010110110",
    "1111011011101000",
    "1111100101000000",
    "1111101110011011",
    "1111110111011000",
    "1111111111011011",
    "1111111001101001",
    "1111110011111110",
    "1111101111011101",
    "1111101011111011",
    "1111101001010011",
    "1111100111100100",
    "1111100110110101",
    "1111100111001100",
    "1111101000100110",
    "1111101010111101",
    "1111101101111110",
    "1111110001010011",
    "1111110100100000",
    "1111110111001010",
    "1111111000111000",
    "1111111001011001",
    "1111111000100100",
    "1111110110100010",
    "1111110011110001",
    "1111110000111100",
    "1111101110110001",
    "1111101101110011",
    "1111101110001010",
    "1111101111100100",
    "1111110001011010",
    "1111110010111100",
    "1111110011011110",
    "1111110010011100",
    "1111101111010111",
    "1111101001111001",
    "1111100001110011",
    "1111010111000110",
    "1111001010001111",
    "1110111100000100",
    "1110101101101000",
    "1110100000000010",
    "1110010100001011",
    "1110001010010011",
    "1110000010001010",
    "1101111011001001",
    "1101110100101001",
    "1101101110001101",
    "1101100111111110",
    "1101100010011100",
    "1101011110010111",
    "1101011100100000",
    "1101011101010100",
    "1101100000111000",
    "1101100110111001",
    "1101101110110011",
    "1101111000000011",
    "1110000010001000",
    "1110001100110011",
    "1110010111111100",
    "1110100011100010",
    "1110101111011111",
    "1110111011101011",
    "1111000111101111",
    "1111010011011010",
    "1111011110011011",
    "1111101000100010",
    "1111110001100101",
    "1111111001011111",
    "1111111111101100",
    "1111111001111111",
    "1111110101001101",
    "1111110001001011",
    "1111101101101100",
    "1111101010101010",
    "1111101000000101",
    "1111100110000001",
    "1111100100101010",
    "1111100100000101",
    "1111100100010010",
    "1111100101010000",
    "1111100110111000",
    "1111101000111100",
    "1111101011010011",
    "1111101101110111",
    "1111110000101001",
    "1111110011101010",
    "1111110111000000",
    "1111111010101101",
    "1111111110111010",
    "1111111100010100",
    "1111110110111110",
    "1111110001001110",
    "1111101011100000",
    "1111100110010101",
    "1111100010010100",
    "1111011111111010",
    "1111011111011001",
    "1111100000110000",
    "1111100011101110",
    "1111100111110111",
    "1111101100101101",
    "1111110001111001",
    "1111110111000101",
    "1111111100000000",
    "1111111111101010",
    "1111111100011001",
    "1111111010100100",
    "1111111010011111",
    "1111111100010100",
    "1111111111111100",
    "1111111010101000",
    "1111110100000010",
    "1111101100100011",
    "1111100100100111",
    "1111011100110101",
    "1111010101110110",
    "1111010000011100",
    "1111001101000100",
    "1111001100000100",
    "1111001101011100",
    "1111010000111001",
    "1111010110000011",
    "1111011100010110",
    "1111100011001010",
    "1111101001110101",
    "1111101111110110",
    "1111110100111011",
    "1111111001000000",
    "1111111100001111",
    "1111111110111011",
    "1111111110101011",
    "1111111100100010",
    "1111111010100011",
    "1111111000101111",
    "1111110111000001",
    "1111110101010011",
    "1111110011100001",
    "1111110001101111",
    "1111110000000100",
    "1111101110101101",
    "1111101101111000",
    "1111101101101100",
    "1111101110001010",
    "1111101111010010",
    "1111110001000011",
    "1111110011011101",
    "1111110110010111",
    "1111111001011111",
    "1111111100010011",
    "1111111110010001",
    "1111111111000000",
    "1111111110010111",
    "1111111100101000",
    "1111111010001110",
    "1111110111100011",
    "1111110100111100",
    "1111110010100011",
    "1111110000011110",
    "1111101110110101",
    "1111101101101100",
    "1111101100111101",
    "1111101100011010",
    "1111101011101011",
    "1111101010100000",
    "1111101000111001",
    "1111100111010000",
    "1111100110010000",
    "1111100110011101",
    "1111101000001100",
    "1111101011011000",
    "1111101111100100",
    "1111110100001001",
    "1111111000011100",
    "1111111100000111",
    "1111111110111111",
    "1111111110111000",
    "1111111101011011",
    "1111111100100000",
    "1111111011111110",
    "1111111011110100",
    "1111111100000010",
    "1111111100101001",
    "1111111101101110",
    "1111111111010000",
    "1111111110110010",
    "1111111100110001",
    "1111111010111110",
    "1111111001110001",
    "1111111001010110",
    "1111111001101000",
    "1111111010010000",
    "1111111010101110",
    "1111111010100010",
    "1111111001011100",
    "1111110111011111",
    "1111110100111111",
    "1111110010010110",
    "1111101111111001",
    "1111101101111001",
    "1111101100100001",
    "1111101011111000",
    "1111101100000011",
    "1111101101001010",
    "1111101111000111",
    "1111110001100110",
    "1111110100000101",
    "1111110101111101",
    "1111110110101100",
    "1111110110000101",
    "1111110100001101",
    "1111110001011100",
    "1111101110001010",
    "1111101010101000",
    "1111100110111011",
    "1111100010110110",
    "1111011101111101",
    "1111010111111001",
    "1111010000011110",
    "1111001000000001",
    "1110111111010010",
    "1110110111001011",
    "1110110000100001",
    "1110101011110111",
    "1110101001001100",
    "1110101000010000",
    "1110101000011101",
    "1110101001011000",
    "1110101010110010",
    "1110101100110011",
    "1110101111101110",
    "1110110011111011",
    "1110111001110000",
    "1111000001011010",
    "1111001010100110",
    "1111010100100101",
    "1111011110001101",
    "1111100110001110",
    "1111101011101110",
    "1111101110001111",
    "1111101110000011",
    "1111101011111111",
    "1111101001001010",
    "1111100110100010",
    "1111100100101100",
    "1111100011101100",
    "1111100011001011",
    "1111100010101011",
    "1111100001110110",
    "1111100000100111",
    "1111011111000100",
    "1111011101010110",
    "1111011011101010",
    "1111011010000100",
    "1111011000101101",
    "1111010111100111",
    "1111010110101101",
    "1111010101111001",
    "1111010100111001",
    "1111010011011010",
    "1111010001010010",
    "1111001110100100",
    "1111001011101000",
    "1111001000111001",
    "1111000110101111",
    "1111000101011000",
    "1111000100110110",
    "1111000101000000",
    "1111000101101110",
    "1111000110110010",
    "1111000111111110",
    "1111001001000001",
    "1111001001101010",
    "1111001001100011",
    "1111001000100101",
    "1111000110110010",
    "1111000100100010",
    "1111000010100010",
    "1111000001101001",
    "1111000010101001",
    "1111000110001001",
    "1111001100010111",
    "1111010101000101",
    "1111011111101100",
    "1111101011011001",
    "1111110111001010",
    "1111111101111100",
    "1111110100110010",
    "1111101101110000",
    "1111101000111000",
    "1111100101110100",
    "1111100011110110",
    "1111100010001011",
    "1111011111111111",
    "1111011100101101",
    "1111011000000011",
    "1111010010000101",
    "1111001011010011",
    "1111000100100000",
    "1110111110101001",
    "1110111010011000",
    "1110110111111010",
    "1110110111000100",
    "1110110111001101",
    "1110110111011111",
    "1110110111010000",
    "1110110110001000",
    "1110110100001010",
    "1110110001100100",
    "1110101110110110",
    "1110101100011001",
    "1110101010100000",
    "1110101001011000",
    "1110101001000001",
    "1110101001011101",
    "1110101010100011",
    "1110101100001110",
    "1110101110010010",
    "1110110000100110",
    "1110110010111001",
    "1110110101000000",
    "1110110110110010",
    "1110111000100000",
    "1110111011011011",
    "1111000010000011",
    "1111001111000010",
    "1111100011101010",
    "1111111110111000",
    "1111100010111000",
    "1111000110011111",
    "1110110000100111",
    "1110100100010010",
    "1110100001011111",
    "1110100101101110",
    "1110101101001010",
    "1110110100010010",
    "1110111000111001",
    "1110111010011110",
    "1110111001100101",
    "1110110111011011",
    "1110110101000011",
    "1110110010111001",
    "1110110001000000",
    "1110101111001101",
    "1110101101011011",
    "1110101011110101",
    "1110101010110100",
    "1110101010100011",
    "1110101010111000",
    "1110101011010011",
    "1110101011011011",
    "1110101011001111",
    "1110101011000010",
    "1110101011001110",
    "1110101100010011",
    "1110101110101001",
    "1110110010101100",
    "1110111000110010",
    "1111000001000101",
    "1111001011001111",
    "1111010110011010",
    "1111100001001111",
    "1111101010000111",
    "1111101111101000",
    "1111110000111111",
    "1111101110010101",
    "1111101000110001",
    "1111100010000000",
    "1111011011111100",
    "1111011000000110",
    "1111010111010011",
    "1111011001100000",
    "1111011101111011",
    "1111100011100110",
    "1111101001100101",
    "1111101111001010",
    "1111110011110011",
    "1111110111001110",
    "1111111001001110",
    "1111111001111011",
    "1111111001101001",
    "1111111000111100",
    "1111111000100001",
    "1111111001000000",
    "1111111010111001",
    "1111111110010100",
    "1111111101000000",
    "1111110111110001",
    "1111110010100111",
    "1111101110001011",
    "1111101010110011",
    "1111101000011101",
    "1111100110111000",
    "1111100101100100",
    "1111100011111100",
    "1111100001101100",
    "1111011110101001",
    "1111011010110101",
    "1111010110101000",
    "1111010010101001",
    "1111001111011100",
    "1111001101100100",
    "1111001101001110",
    "1111001110001111",
    "1111010000001100",
    "1111010010011100",
    "1111010100011100",
    "1111010101101010",
    "1111010101110001",
    "1111010100011101",
    "1111010001100010",
    "1111001100111000",
    "1111000110100111",
    "1110111111001100",
    "1110110111001110",
    "1110101111100100",
    "1110101000111110",
    "1110100011110110",
    "1110100000001111",
    "1110011101110111",
    "1110011100010011",
    "1110011011000110",
    "1110011001111111",
    "1110011000111110",
    "1110011000001011",
    "1110010111111110",
    "1110011000101100",
    "1110011010101011",
    "1110011110000000",
    "1110100010100010",
    "1110100111101111",
    "1110101101000000",
    "1110110001110110",
    "1110110110000000",
    "1110111001011110",
    "1110111100011100",
    "1110111111000000",
    "1111000001001000",
    "1111000010100111",
    "1111000011010101",
    "1111000011001111",
    "1111000010100001",
    "1111000001100001",
    "1111000000100100",
    "1110111111111011",
    "1110111111101000",
    "1110111111101110",
    "1111000000010100",
    "1111000001100110",
    "1111000011101111",
    "1111000110111011",
    "1111001011000110",
    "1111010000000010",
    "1111010101011101",
    "1111011011000001",
    "1111100000010111",
    "1111100101001101",
    "1111101001001100",
    "1111101011111000",
    "1111101100101101",
    "1111101011001101",
    "1111100111001100",
    "1111100000110110",
    "1111011000110000",
    "1111001111110101",
    "1111000111000011",
    "1110111111010100",
    "1110111001011000",
    "1110110101100101",
    "1110110100000110",
    "1110110100110110",
    "1110110111101000",
    "1110111100001111",
    "1111000010010111",
    "1111001001100111",
    "1111010001100110",
    "1111011001110100",
    "1111100001110000",
    "1111101000110110",
    "1111101110100010",
    "1111110010010110",
    "1111110011111101",
    "1111110011010101",
    "1111110000101110",
    "1111101100101000",
    "1111100111101110",
    "1111100010110011",
    "1111011110100100",
    "1111011011100011",
    "1111011010001011",
    "1111011010100101",
    "1111011100110000",
    "1111100000010100",
    "1111100100101110",
    "1111101001010010",
    "1111101101011011",
    "1111110000101111",
    "1111110011000111",
    "1111110100101110",
    "1111110101111010",
    "1111110110111101",
    "1111111000000010",
    "1111111001001001",
    "1111111010000010",
    "1111111010100001",
    "1111111010100000",
    "1111111010000000",
    "1111111001010000",
    "1111111000011011",
    "1111110111101000",
    "1111110110110100",
    "1111110101111000",
    "1111110100101011",
    "1111110011010010",
    "1111110001111111",
    "1111110001010100",
    "1111110001110000",
    "1111110011101011",
    "1111110111001000",
    "1111111011110011",
    "1111111110110110",
    "1111111001011111",
    "1111110100100001",
    "1111110000001000",
    "1111101100001101",
    "1111101000101000",
    "1111100101010101",
    "1111100010010010",
    "1111011111100001",
    "1111011100111100",
    "1111011010010001",
    "1111010111001110",
    "1111010011100010",
    "1111001111001111",
    "1111001010100110",
    "1111000110001000",
    "1111000010100001",
    "1111000000010111",
    "1111000000001111",
    "1111000010100001",
    "1111000111010011",
    "1111001110011001",
    "1111010111001110",
    "1111100000110110",
    "1111101010010001",
    "1111110010100000",
    "1111111000111011",
    "1111111101011011",
    "1111111111100111",
    "1111111101100111",
    "1111111011111000",
    "1111111001111111",
    "1111110111110110",
    "1111110101101110",
    "1111110100000011",
    "1111110011001100",
    "1111110011010110",
    "1111110100010111",
    "1111110101110111",
    "1111110111010111",
    "1111111000100001",
    "1111111001001110",
    "1111111001111100",
    "1111111011100110",
    "1111111111011101",
    "1111111001100000",
    "1111101111000011",
    "1111100001101110",
    "1111010010111001",
    "1111000100010101",
    "1110110111110010",
    "1110101110011111",
    "1110101000111010",
    "1110100110101100",
    "1110100110111111",
    "1110101000111010",
    "1110101011101000",
    "1110101110101110",
    "1110110010001010",
    "1110110110000001",
    "1110111010011011",
    "1110111111010111",
    "1111000100100010",
    "1111001001100010",
    "1111001110000000",
    "1111010001101110",
    "1111010100011101",
    "1111010110000011",
    "1111010110010010",
    "1111010100111011",
    "1111010001110001",
    "1111001100110101",
    "1111000110001001",
    "1110111110000101",
    "1110110101001000",
    "1110101011110111",
    "1110100010111011",
    "1110011010111010",
    "1110010100010101",
    "1110001111110000",
    "1110001101100001",
    "1110001101111000",
    "1110010000101110",
    "1110010101101110",
    "1110011100011011",
    "1110100100011100",
    "1110101101011001",
    "1110110110111100",
    "1111000000100110",
    "1111001001101101",
    "1111010001100111",
    "1111010111111001",
    "1111011100011001",
    "1111011111100100",
    "1111100010000101",
    "1111100100101001",
    "1111100111101010",
    "1111101011001111",
    "1111101111000111",
    "1111110011000001",
    "1111110110101001",
    "1111111001110011",
    "1111111100010111",
    "1111111110001010",
    "1111111110111011",
    "1111111110001101",
    "1111111011100110",
    "1111110110101110",
    "1111101111011111",
    "1111100110001011",
    "1111011011100001",
    "1111010000011110",
    "1111000110001000",
    "1110111101100001",
    "1110110111010110",
    "1110110011111001",
    "1110110010110011",
    "1110110011010111",
    "1110110100100111",
    "1110110101110001",
    "1110110110010110",
    "1110110110010000",
    "1110110101101111",
    "1110110101000110",
    "1110110100101111",
    "1110110101000000",
    "1110110110001000",
    "1110111000100000",
    "1110111100011110",
    "1111000010010100",
    "1111001010000111",
    "1111010011110001",
    "1111011110110110",
    "1111101010110001",
    "1111110110110100",
    "1111111101100101",
    "1111110011000101",
    "1111101001111111",
    "1111100010011111",
    "1111011100100110",
    "1111011000010110",
    "1111010101101001",
    "1111010100010010",
    "1111010100000011",
    "1111010100100111",
    "1111010101100010",
    "1111010110011101",
    "1111010110111011",
    "1111010110101000",
    "1111010101011000",
    "1111010011001010",
    "1111010000000111",
    "1111001100100001",
    "1111001000110010",
    "1111000101010010",
    "1111000010001101",
    "1110111111101100",
    "1110111101101011",
    "1110111011111010",
    "1110111010000110",
    "1110110111111110",
    "1110110101011111",
    "1110110010101011",
    "1110101111110001",
    "1110101101000111",
    "1110101010110101",
    "1110101001000001",
    "1110100111100011",
    "1110100110010000",
    "1110100100111011",
    "1110100011011111",
    "1110100010000010",
    "1110100000101011",
    "1110011111100100",
    "1110011110111010",
    "1110011110101011",
    "1110011110111010",
    "1110011111100110",
    "1110100000101110",
    "1110100010011010",
    "1110100100110011",
    "1110101000001100",
    "1110101101011011",
    "1110110101110111",
    "1111000011001000",
    "1111010101111011",
    "1111101101101011",
    "1111110111100111",
    "1111011101001001",
    "1111000110001110",
    "1110110101011000",
    "1110101011011000",
    "1110100111001110",
    "1110100110111001",
    "1110101000011000",
    "1110101010001110",
    "1110101011111000",
    "1110101101011110",
    "1110101111010110",
    "1110110001110000",
    "1110110100011101",
    "1110110111000001",
    "1110111000111010",
    "1110111001111010",
    "1110111010001111",
    "1110111010010011",
    "1110111010100010",
    "1110111011000110",
    "1110111011111010",
    "1110111100110101",
    "1110111101101101",
    "1110111110100011",
    "1110111111010111",
    "1111000000010101",
    "1111000001101011",
    "1111000011011111",
    "1111000110000100",
    "1111001001100111",
    "1111001110001001",
    "1111010011010111",
    "1111011000101100",
    "1111011101010010",
    "1111100000010101",
    "1111100001010100",
    "1111100000000111",
    "1111011101001001",
    "1111011001001110",
    "1111010101010111",
    "1111010010011100",
    "1111010001000000",
    "1111010001001100",
    "1111010010101110",
    "1111010101010010",
    "1111011000100111",
    "1111011100100011",
    "1111100001000111",
    "1111100110010000",
    "1111101011111011",
    "1111110010000010",
    "1111111000011010",
    "1111111110111100",
    "1111111010100010",
    "1111110100001101",
    "1111101110010011",
    "1111101001000010",
    "1111100100110011",
    "1111100001110100",
    "1111100000010101",
    "1111100000011001",
    "1111100001111000",
    "1111100100100111",
    "1111101000001001",
    "1111101100000000",
    "1111101111101001",
    "1111110010101010",
    "1111110100110010",
    "1111110101111010",
    "1111110110001010",
    "1111110101110001",
    "1111110101000000",
    "1111110100001001",
    "1111110011010010",
    "1111110010100010",
    "1111110001110100",
    "1111110001000010",
    "1111101111111110",
    "1111101110010101",
    "1111101011110100",
    "1111101000000010",
    "1111100010100111",
    "1111011011011000",
    "1111010010010000",
    "1111000111100010",
    "1110111011101011",
    "1110101111010001",
    "1110100011000000",
    "1110010111100010",
    "1110001101010010",
    "1110000100011100",
    "1101111100110101",
    "1101110110010000",
    "1101110000011111",
    "1101101011011011",
    "1101100111001110",
    "1101100100001110",
    "1101100010111000",
    "1101100011100100",
    "1101100110100100",
    "1101101011101111",
    "1101110010100110",
    "1101111010011011",
    "1110000010010111",
    "1110001001110000",
    "1110010000010010",
    "1110010110001011",
    "1110011011111101",
    "1110100010010000",
    "1110101001100000",
    "1110110001101110",
    "1110111010101101",
    "1111000100001011",
    "1111001101110111",
    "1111010111110001",
    "1111100001111001",
    "1111101100001011",
    "1111110110010101",
    "1111111111110111",
    "1111110111101111",
    "1111110000111100",
    "1111101011110100",
    "1111101000001011",
    "1111100101101100",
    "1111100100001011",
    "1111100011100110",
    "1111100100001011",
    "1111100110001011",
    "1111101001110101",
    "1111101111000110",
    "1111110101101010",
    "1111111100111010",
    "1111111011110011",
    "1111110101010010",
    "1111110000000111",
    "1111101100100111",
    "1111101010111001",
    "1111101010110100",
    "1111101100000010",
    "1111101110001000",
    "1111110000101110",
    "1111110011011100",
    "1111110101111110",
    "1111111000001000",
    "1111111001110010",
    "1111111010111011",
    "1111111011101000",
    "1111111100000000",
    "1111111100001001",
    "1111111100001001",
    "1111111100000000",
    "1111111011101101",
    "1111111011001001",
    "1111111010001101",
    "1111111000101011",
    "1111110110010100",
    "1111110010111101",
    "1111101110011110",
    "1111101000111111",
    "1111100010111001",
    "1111011100110101",
    "1111010111100010",
    "1111010011101110",
    "1111010001110011",
    "1111010001111110",
    "1111010100000000",
    "1111010111011111",
    "1111011011110010",
    "1111100000010100",
    "1111100100011111",
    "1111100111111100",
    "1111101010100111",
    "1111101100110010",
    "1111101110111100",
    "1111110001101000",
    "1111110101001010",
    "1111111001100001",
    "1111111110010111",
    "1111111100110010",
    "1111111000100011",
    "1111110101001100",
    "1111110010111010",
    "1111110001101111",
    "1111110001101010",
    "1111110010101001",
    "1111110100100000",
    "1111110110111011",
    "1111111001011111",
    "1111111011100111",
    "1111111100111001",
    "1111111101000111",
    "1111111100010001",
    "1111111010101010",
    "1111111000100100",
    "1111110110010000",
    "1111110011111010",
    "1111110001110000",
    "1111101111111100",
    "1111101110101110",
    "1111101110001110",
    "1111101110011111",
    "1111101111010000",
    "1111110000001011",
    "1111110000111011",
    "1111110001010000",
    "1111110001000110",
    "1111110000011100",
    "1111101111010111",
    "1111101101110111",
    "1111101100000110",
    "1111101010010111",
    "1111101001001001",
    "1111101000111110",
    "1111101010001110",
    "1111101101000000",
    "1111110000111111",
    "1111110101100101",
    "1111111010000011",
    "1111111101110010",
    "1111111111100001",
    "1111111101111100",
    "1111111101010001",
    "1111111101000101",
    "1111111101000111",
    "1111111101001011",
    "1111111101010001",
    "1111111101100100",
    "1111111110001110",
    "1111111111011110",
    "1111111110101010",
    "1111111100010101",
    "1111111001101111",
    "1111110111010000",
    "1111110101010010",
    "1111110100000011",
    "1111110011100001",
    "1111110011100010",
    "1111110011101110",
    "1111110011110011",
    "1111110011101100",
    "1111110011011101",
    "1111110011011011",
    "1111110011111001",
    "1111110101000100",
    "1111110110111111",
    "1111111001011100",
    "1111111100000011",
    "1111111110011101",
    "1111111111101100",
    "1111111110101010",
    "1111111110100010",
    "1111111111001111",
    "1111111111010001",
    "1111111101001010",
    "1111111010011000",
    "1111110110110101",
    "1111110010100011",
    "1111101101011011",
    "1111100111100001",
    "1111100000110101",
    "1111011001011110",
    "1111010001110001",
    "1111001010000010",
    "1111000010110011",
    "1110111100011011",
    "1110110111010011",
    "1110110011101001",
    "1110110001011001",
    "1110110000001111",
    "1110101111110000",
    "1110101111010111",
    "1110101110111000",
    "1110101110010010",
    "1110101101111101",
    "1110101110011110",
    "1110110000100011",
    "1110110100100111",
    "1110111010110100",
    "1111000010111000",
    "1111001100000101",
    "1111010101011101",
    "1111011101111101",
    "1111100100101001",
    "1111101000111111",
    "1111101010111101",
    "1111101010110111",
    "1111101001011010",
    "1111100111010000",
    "1111100100111001",
    "1111100010100010",
    "1111100000001101",
    "1111011101110011",
    "1111011011010100",
    "1111011000110010",
    "1111010110100000",
    "1111010100110001",
    "1111010011110100",
    "1111010011110001",
    "1111010100100000",
    "1111010101101111",
    "1111010111000100",
    "1111011000000011",
    "1111011000001001",
    "1111010110111110",
    "1111010100001101",
    "1111001111110110",
    "1111001010010001",
    "1111000100000000",
    "1110111101110011",
    "1110111000010110",
    "1110110100001000",
    "1110110001011010",
    "1110110000010100",
    "1110110000110011",
    "1110110010110100",
    "1110110110010010",
    "1110111010111010",
    "1111000000011001",
    "1111000110001001",
    "1111001011100101",
    "1111010000000000",
    "1111010010111110",
    "1111010100001110",
    "1111010011111000",
    "1111010010010100",
    "1111010000010010",
    "1111001110100110",
    "1111001110000100",
    "1111001111010110",
    "1111010010111001",
    "1111011000110101",
    "1111100001000000",
    "1111101010110011",
    "1111110101010110",
    "1111111111101000",
    "1111110111001011",
    "1111101111101101",
    "1111101010000100",
    "1111100101111011",
    "1111100010101001",
    "1111011111100001",
    "1111011011111111",
    "1111010111101101",
    "1111010010101110",
    "1111001101001111",
    "1111000111110101",
    "1111000011000000",
    "1110111111010010",
    "1110111100111000",
    "1110111011110011",
    "1110111011101101",
    "1110111100000010",
    "1110111100001010",
    "1110111011100101",
    "1110111010000001",
    "1110110111011010",
    "1110110100000011",
    "1110110000011001",
    "1110101100111101",
    "1110101010001110",
    "1110101000011101",
    "1110100111110100",
    "1110101000010001",
    "1110101001101011",
    "1110101011110010",
    "1110101110010100",
    "1110110001000000",
    "1110110011100111",
    "1110110110000110",
    "1110111000100111",
    "1110111100001010",
    "1111000010101100",
    "1111001110001010",
    "1111011111100110",
    "1111110110011100",
    "1111101111101011",
    "1111010110011010",
    "1111000001010101",
    "1110110011000011",
    "1110101100000001",
    "1110101010111000",
    "1110101101010001",
    "1110110000101110",
    "1110110011100010",
    "1110110101000011",
    "1110110101010111",
    "1110110100111001",
    "1110110100001011",
    "1110110011010011",
    "1110110010010000",
    "1110110000111110",
    "1110101111100011",
    "1110101110001111",
    "1110101101011001",
    "1110101101010001",
    "1110101101101110",
    "1110101110011110",
    "1110101111001000",
    "1110101111101000",
    "1110101111111101",
    "1110110000010100",
    "1110110000111001",
    "1110110001111110",
    "1110110011101010",
    "1110110110001101",
    "1110111001101101",
    "1110111110010110",
    "1111000100001011",
    "1111001011001001",
    "1111010010110110",
    "1111011010101101",
    "1111100001110001",
    "1111100111001011",
    "1111101010010001",
    "1111101010111001",
    "1111101001011111",
    "1111100110110101",
    "1111100011111011",
    "1111100001100001",
    "1111100000000111",
    "1111011111111011",
    "1111100000111001",
    "1111100010110100",
    "1111100101011101",
    "1111101000011110",
    "1111101011100111",
    "1111101110110001",
    "1111110001111100",
    "1111110101010000",
    "1111111000111000",
    "1111111101000001",
    "1111111110001110",
    "1111111001001000",
    "1111110100000000",
    "1111101111011000",
    "1111101011110000",
    "1111101001010110",
    "1111101000001101",
    "1111101000000010",
    "1111101000011010",
    "1111101000110000",
    "1111101000101001",
    "1111100111110010",
    "1111100110000011",
    "1111100011100111",
    "1111100000101110",
    "1111011101101101",
    "1111011010110111",
    "1111011000010110",
    "1111010110001110",
    "1111010100100010",
    "1111010011001111",
    "1111010010001111",
    "1111010001010111",
    "1111010000010100",
    "1111001110101110",
    "1111001100001100",
    "1111001000010110",
    "1111000011000011",
    "1110111100011001",
    "1110110100101010",
    "1110101100011001",
    "1110100100001101",
    "1110011100110111",
    "1110010111000011",
    "1110010011001111",
    "1110010001100111",
    "1110010010000110",
    "1110010100010101",
    "1110010111110010",
    "1110011100000010",
    "1110100000110000",
    "1110100101101001",
    "1110101010100011",
    "1110101111000111",
    "1110110010110110",
    "1110110101010000",
    "1110110101111110",
    "1110110100111011",
    "1110110010100010",
    "1110101111011010",
    "1110101100001111",
    "1110101001011101",
    "1110100111010101",
    "1110100110000100",
    "1110100101111011",
    "1110100111001101",
    "1110101010010001",
    "1110101111001101",
    "1110110101110110",
    "1110111101100100",
    "1111000101100111",
    "1111001101001001",
    "1111010011011111",
    "1111011000010000",
    "1111011011001110",
    "1111011100100001",
    "1111011100011011",
    "1111011011010100",
    "1111011001101101",
    "1111011000000001",
    "1111010110100111",
    "1111010101100101",
    "1111010100101111",
    "1111010011101111",
    "1111010010001011",
    "1111001111110101",
    "1111001100101000",
    "1111001000111010",
    "1111000101001101",
    "1111000001111101",
    "1110111111100100",
    "1110111110010100",
    "1110111110001010",
    "1110111111000101",
    "1111000000111110",
    "1111000011101010",
    "1111000111000011",
    "1111001010111100",
    "1111001111001101",
    "1111010011101111",
    "1111011000010000",
    "1111011100011001",
    "1111011111110011",
    "1111100010000110",
    "1111100011000011",
    "1111100010100111",
    "1111100001000010",
    "1111011110110000",
    "1111011100010111",
    "1111011010010110",
    "1111011000111111",
    "1111011000011010",
    "1111011000100010",
    "1111011001010001",
    "1111011010100000",
    "1111011100000111",
    "1111011110000000",
    "1111100000000111",
    "1111100010010100",
    "1111100100011101",
    "1111100110101000",
    "1111101001000001",
    "1111101011111100",
    "1111101111101111",
    "1111110100011001",
    "1111111001100011",
    "1111111110011111",
    "1111111101100111",
    "1111111011100010",
    "1111111011100110",
    "1111111101101110",
    "1111111110100011",
    "1111111001111111",
    "1111110101010001",
    "1111110000111101",
    "1111101101011100",
    "1111101010111100",
    "1111101001100000",
    "1111101001001010",
    "1111101001110010",
    "1111101011010011",
    "1111101101100101",
    "1111110000011100",
    "1111110011110000",
    "1111110111011001",
    "1111111011010010",
    "1111111111010110",
    "1111111100011010",
    "1111111000001001",
    "1111110011111100",
    "1111101111111000",
    "1111101011111101",
    "1111101000000101",
    "1111100100000000",
    "1111011111011110",
    "1111011010001100",
    "1111010100001110",
    "1111001101110010",
    "1111000111010001",
    "1111000001010111",
    "1110111100100101",
    "1110111001011101",
    "1110111000011000",
    "1110111001101000",
    "1110111101010110",
    "1111000011011101",
    "1111001011101111",
    "1111010101100100",
    "1111100000000101",
    "1111101010010011",
    "1111110011010101",
    "1111111010100100",
    "1111111111110110",
    "1111111100100001",
    "1111111010001101",
    "1111111000100101",
    "1111110111010100",
    "1111110110010001",
    "1111110101011111",
    "1111110101001011",
    "1111110101011011",
    "1111110110001010",
    "1111110111000101",
    "1111110111111001",
    "1111111000010010",
    "1111111000001111",
    "1111111000001011",
    "1111111000111100",
    "1111111011100000",
    "1111111111011010",
    "1111110111110000",
    "1111101110001101",
    "1111100100000101",
    "1111011010110010",
    "1111010011101001",
    "1111001111001010",
    "1111001101010010",
    "1111001101010010",
    "1111001110010010",
    "1111001111011111",
    "1111010000010111",
    "1111010000110001",
    "1111010000110000",
    "1111010000100001",
    "1111010000001101",
    "1111001111111011",
    "1111001111101110",
    "1111001111011111",
    "1111001111010001",
    "1111001110111011",
    "1111001110011100",
    "1111001101100110",
    "1111001100001001",
    "1111001001110100",
    "1111000110011101",
    "1111000010000011",
    "1110111100100110",
    "1110110110001011",
    "1110101110110110",
    "1110100110110010",
    "1110011110010111",
    "1110010110001011",
    "1110001110111010",
    "1110001001010110",
    "1110000101111110",
    "1110000101000001",
    "1110000110100101",
    "1110001010100000",
    "1110010000101100",
    "1110011000111010",
    "1110100010110001",
    "1110101101100001",
    "1110111000010110",
    "1111000010010101",
    "1111001010110000",
    "1111010001010000",
    "1111010101111011",
    "1111011001000010",
    "1111011011000100",
    "1111011100011100",
    "1111011101101001",
    "1111011111000111",
    "1111100001001010",
    "1111100100001010",
    "1111101000000101",
    "1111101100110001",
    "1111110001101010",
    "1111110110001010",
    "1111111001100011",
    "1111111011010101",
    "1111111011001001",
    "1111111000101111",
    "1111110011111101",
    "1111101100101101",
    "1111100011001011",
    "1111010111110111",
    "1111001011101101",
    "1110111111111011",
    "1110110101101010",
    "1110101101110011",
    "1110101000101101",
    "1110100110001001",
    "1110100101100100",
    "1110100110000110",
    "1110100111000011",
    "1110100111110111",
    "1110101000010011",
    "1110101000011011",
    "1110101000011110",
    "1110101000111010",
    "1110101010000001",
    "1110101100000111",
    "1110101111010111",
    "1110110011110011",
    "1110111001100000",
    "1111000000011111",
    "1111001000110000",
    "1111010010001000",
    "1111011100010100",
    "1111100110111111",
    "1111110001110011",
    "1111111100100001",
    "1111111000111111",
    "1111101110111101",
    "1111100101100010",
    "1111011101000111",
    "1111010110001000",
    "1111010000111110",
    "1111001101111010",
    "1111001100110111",
    "1111001101011100",
    "1111001111000111",
    "1111010001010010",
    "1111010011011111",
    "1111010101011000",
    "1111010110110001",
    "1111010111100000",
    "1111010111100000",
    "1111010110101010",
    "1111010100111011",
    "1111010010010101",
    "1111001111000000",
    "1111001011000111",
    "1111000110110010",
    "1111000010001010",
    "1110111101010010",
    "1110111000001110",
    "1110110011001111",
    "1110101110100100",
    "1110101010101011",
    "1110100111110101",
    "1110100110001000",
    "1110100101011010",
    "1110100101010101",
    "1110100101100000",
    "1110100101100111",
    "1110100101011111",
    "1110100101001001",
    "1110100100101111",
    "1110100100011010",
    "1110100100001110",
    "1110100100001110",
    "1110100100010011",
    "1110100100011010",
    "1110100100100111",
    "1110100101001000",
    "1110100110001011",
    "1110101000001011",
    "1110101011100101",
    "1110110001011100",
    "1110111011010011",
    "1111001010011101",
    "1111011111010010",
    "1111111000101000",
    "1111101011111100",
    "1111010001111001",
    "1110111100100011",
    "1110101110000000",
    "1110100110100111",
    "1110100100111001",
    "1110100110101010",
    "1110101001101111",
    "1110101100110000",
    "1110101111010100",
    "1110110001101001",
    "1110110100001101",
    "1110110111001101",
    "1110111010010110",
    "1110111101000100",
    "1110111110110011",
    "1110111111010001",
    "1110111110101001",
    "1110111101011110",
    "1110111100001111",
    "1110111011001110",
    "1110111010011101",
    "1110111001111100",
    "1110111001101011",
    "1110111001101111",
    "1110111010001011",
    "1110111011001110",
    "1110111101001110",
    "1111000000011100",
    "1111000101000000",
    "1111001010101000",
    "1111010000100110",
    "1111010110000011",
    "1111011001111100",
    "1111011011100110",
    "1111011010101010",
    "1111010111011011",
    "1111010010101011",
    "1111001101011001",
    "1111001000101111",
    "1111000101101010",
    "1111000100110100",
    "1111000110011011",
    "1111001010010100",
    "1111001111111111",
    "1111010110110110",
    "1111011110011011",
    "1111100110010101",
    "1111101110010001",
    "1111110101111100",
    "1111111101000110",
    "1111111100100000",
    "1111110111000110",
    "1111110010101100",
    "1111101111001011",
    "1111101100010100",
    "1111101001110001",
    "1111100111011010",
    "1111100101011000",
    "1111100100000011",
    "1111100011111000",
    "1111100101001001",
    "1111100111111111",
    "1111101100000011",
    "1111110000101111",
    "1111110101010010",
    "1111111001000001",
    "1111111011011101",
    "1111111100011001",
    "1111111011111010",
    "1111111010010100",
    "1111111000000011",
    "1111110101100010",
    "1111110011000100",
    "1111110000101101",
    "1111101110010000",
    "1111101011011001",
    "1111100111110100",
    "1111100011010011",
    "1111011101110111",
    "1111010111101100",
    "1111010001000011",
    "1111001010011000",
    "1111000011110110",
    "1110111101101001",
    "1110110111110111",
    "1110110010011101",
    "1110101101010110",
    "1110101000010101",
    "1110100011000011",
    "1110011101001100",
    "1110010110011011",
    "1110001110101001",
    "1110000101111110",
    "1101111100110011",
    "1101110011110100",
    "1101101011110011",
    "1101100101100010",
    "1101100001100110",
    "1101100000010001",
    "1101100001100001",
    "1101100100111110",
    "1101101010001001",
    "1101110000011100",
    "1101110111100010",
    "1101111111010010",
    "1110000111101101",
    "1110010000111011",
    "1110011010111100",
    "1110100101101100",
    "1110110001000010",
    "1110111100101101",
    "1111001000011110",
    "1111010100001011",
    "1111011111011010",
    "1111101001101101",
    "1111110010100001",
    "1111111001010101",
    "1111111101111000",
    "1111111111101010",
    "1111111110111101",
    "1111111111001111",
    "1111111111110000",
    "1111111111111101",
    "1111111111101100",
    "1111111111000101",
    "1111111110011100",
    "1111111110000011",
    "1111111110000110",
    "1111111110100100",
    "1111111111010110",
    "1111111111101011",
    "1111111110101001",
    "1111111101100010",
    "1111111100010010",
    "1111111010110101",
    "1111111001001101",
    "1111110111100111",
    "1111110110010001",
    "1111110101011100",
    "1111110101011001",
    "1111110110001010",
    "1111110111101000",
    "1111111001100101",
    "1111111011101100",
    "1111111101101010",
    "1111111111001011",
    "1111111111111110",
    "1111111111110101",
    "1111111110100001",
    "1111111011111111",
    "1111111000010011",
    "1111110011101011",
    "1111101110011011",
    "1111101000111100",
    "1111100011101110",
    "1111011111000101",
    "1111011011011000",
    "1111011000101101",
    "1111010111001001",
    "1111010110100100",
    "1111010110111011",
    "1111011000001100",
    "1111011010010110",
    "1111011101010010",
    "1111100000101110",
    "1111100100001110",
    "1111100111010111",
    "1111101001110100",
    "1111101011100110",
    "1111101100111101",
    "1111101110001011",
    "1111101111100010",
    "1111110001000100",
    "1111110010101110",
    "1111110100011110",
    "1111110110010111",
    "1111111000100011",
    "1111111011000111",
    "1111111101111101",
    "1111111111001010",
    "1111111100110101",
    "1111111011011001",
    "1111111010111111",
    "1111111011100001",
    "1111111100101011",
    "1111111110000011",
    "1111111111010011",
    "1111111111110110",
    "1111111111101101",
    "1111111111100010",
    "1111111101111001",
    "1111111011011100",
    "1111111000011011",
    "1111110101010000",
    "1111110010010100",
    "1111101111111001",
    "1111101110000111",
    "1111101100111100",
    "1111101100010000",
    "1111101011111100",
    "1111101011110101",
    "1111101011101101",
    "1111101011010100",
    "1111101010100100",
    "1111101001100000",
    "1111101000011010",
    "1111100111110010",
    "1111101000001101",
    "1111101010000110",
    "1111101101100100",
    "1111110010010111",
    "1111110111110110",
    "1111111101010100",
    "1111111101110110",
    "1111111010001101",
    "1111110111111010",
    "1111110110111101",
    "1111110111001101",
    "1111111000011001",
    "1111111010010100",
    "1111111100110100",
    "1111111111110001",
    "1111111100110111",
    "1111111001010110",
    "1111110101110101",
    "1111110010100111",
    "1111110000000000",
    "1111101110010000",
    "1111101101100001",
    "1111101101110101",
    "1111101111001011",
    "1111110001011011",
    "1111110100010111",
    "1111110111101111",
    "1111111011010001",
    "1111111110100010",
    "1111111110101111",
    "1111111100110101",
    "1111111011110010",
    "1111111011100011",
    "1111111011110110",
    "1111111100011001",
    "1111111100111100",
    "1111111101010000",
    "1111111101010010",
    "1111111101000100",
    "1111111100100111",
    "1111111100000011",
    "1111111011011110",
    "1111111011000111",
    "1111111011001100",
    "1111111100000011",
    "1111111110000010",
    "1111111110100010",
    "1111111001100000",
    "1111110010110110",
    "1111101010101100",
    "1111100001010100",
    "1111010111000011",
    "1111001100011110",
    "1111000010010111",
    "1110111001100011",
    "1110110010101110",
    "1110101110011001",
    "1110101100101011",
    "1110101101001100",
    "1110101111001100",
    "1110110001101011",
    "1110110011101110",
    "1110110100111011",
    "1110110101011000",
    "1110110101101100",
    "1110110110110001",
    "1110111001010101",
    "1110111101101110",
    "1111000011110100",
    "1111001010111000",
    "1111010010000101",
    "1111011000100101",
    "1111011101110010",
    "1111100001100010",
    "1111100011111011",
    "1111100101001101",
    "1111100101101111",
    "1111100101101111",
    "1111100101010011",
    "1111100100010011",
    "1111100010101110",
    "1111100000011111",
    "1111011101110111",
    "1111011011000100",
    "1111011000011000",
    "1111010101110110",
    "1111010011011010",
    "1111010000110110",
    "1111001110000111",
    "1111001011001111",
    "1111001000100111",
    "1111000110100100",
    "1111000101010010",
    "1111000100101010",
    "1111000100010010",
    "1111000011100001",
    "1111000001110011",
    "1110111110110101",
    "1110111010101011",
    "1110110101110010",
    "1110110000101100",
    "1110101011111010",
    "1110100111110100",
    "1110100100101010",
    "1110100010101001",
    "1110100001110110",
    "1110100010100001",
    "1110100100110111",
    "1110101001000111",
    "1110101111010111",
    "1110110111100000",
    "1111000001000111",
    "1111001011010100",
    "1111010101001101",
    "1111011101101110",
    "1111100100010010",
    "1111101000101100",
    "1111101011010101",
    "1111101100111101",
    "1111101110010110",
    "1111110000000010",
    "1111110010001000",
    "1111110100010111",
    "1111110110010011",
    "1111110111101001",
    "1111111000011101",
    "1111111001001101",
    "1111111010100000",
    "1111111100111110",
    "1111111110111111",
    "1111111001011011",
    "1111110010100111",
    "1111101011000000",
    "1111100011000001",
    "1111011011000010",
    "1111010011010011",
    "1111001100001001",
    "1111000101111001",
    "1111000000111101",
    "1110111101101011",
    "1110111100010001",
    "1110111100100011",
    "1110111110000000",
    "1110111111111011",
    "1111000001100010",
    "1111000010001101",
    "1111000001100111",
    "1110111111110101",
    "1110111101000100",
    "1110111001110010",
    "1110110110010110",
    "1110110011001010",
    "1110110000011110",
    "1110101110010111",
    "1110101100111101",
    "1110101100001110",
    "1110101100000111",
    "1110101100100110",
    "1110101101101101",
    "1110101111011010",
    "1110110001111000",
    "1110110101001101",
    "1110111010001001",
    "1111000010001010",
    "1111001110110001",
    "1111100000101001",
    "1111110111000110",
    "1111110000000100",
    "1111011000000100",
    "1111000100001011",
    "1110110110100101",
    "1110101111110000",
    "1110101110001100",
    "1110101111101100",
    "1110110010000010",
    "1110110011110001",
    "1110110100011111",
    "1110110100011000",
    "1110110100000001",
    "1110110011101111",
    "1110110011011101",
    "1110110010111001",
    "1110110001110100",
    "1110110000001111",
    "1110101110011110",
    "1110101101000010",
    "1110101100001111",
    "1110101100001001",
    "1110101100011100",
    "1110101100111010",
    "1110101101010111",
    "1110101101111011",
    "1110101110101101",
    "1110101111110101",
    "1110110001011100",
    "1110110011011111",
    "1110110101111110",
    "1110111000110100",
    "1110111100001001",
    "1111000000000101",
    "1111000100110100",
    "1111001010001100",
    "1111001111101110",
    "1111010100101100",
    "1111011000010011",
    "1111011010000110",
    "1111011010000001",
    "1111011000101100",
    "1111010110111111",
    "1111010101110111",
    "1111010101111100",
    "1111010111011010",
    "1111011010000001",
    "1111011101011100",
    "1111100001010100",
    "1111100101010101",
    "1111101001011011",
    "1111101101100100",
    "1111110001110110",
    "1111110110010100",
    "1111111011000000",
    "1111111111110101",
    "1111111011010011",
    "1111110110100110",
    "1111110010010001",
    "1111101110101001",
    "1111101100000110",
    "1111101010111101",
    "1111101011010101",
    "1111101101000110",
    "1111101111110100",
    "1111110010110100",
    "1111110101010100",
    "1111110110101011",
    "1111110110011010",
    "1111110100010001",
    "1111110000010010",
    "1111101010101010",
    "1111100011110001",
    "1111011100001001",
    "1111010100010101",
    "1111001100111010",
    "1111000110011101",
    "1111000001010100",
    "1110111101110011",
    "1110111011111101",
    "1110111011101011",
    "1110111100100001",
    "1110111101110011",
    "1110111110101110",
    "1110111110100001",
    "1110111100101110",
    "1110111001011000",
    "1110110100110110",
    "1110101111111101",
    "1110101011011110",
    "1110100111111100",
    "1110100101100010",
    "1110100100000011",
    "1110100011001011",
    "1110100010100111",
    "1110100010001010",
    "1110100001101100",
    "1110100001001101",
    "1110100000101011",
    "1110100000000111",
    "1110011111100011",
    "1110011111001000",
    "1110011111000100",
    "1110011111011111",
    "1110100000100001",
    "1110100010001101",
    "1110100100100100",
    "1110100111101000",
    "1110101011011001",
    "1110101111110101",
    "1110110100101100",
    "1110111001101010",
    "1110111110010111",
    "1111000010010111",
    "1111000101011101",
    "1111000111100011",
    "1111001000110100",
    "1111001001100011",
    "1111001010000001",
    "1111001010100101",
    "1111001011011000",
    "1111001100100110",
    "1111001110001101",
    "1111010000000010",
    "1111010001101100",
    "1111010010110001",
    "1111010010110100",
    "1111010001100100",
    "1111001110111011",
    "1111001011001010",
    "1111000110101111",
    "1111000010010000",
    "1110111110010100",
    "1110111011011101",
    "1110111001111010",
    "1110111001110000",
    "1110111010111000",
    "1110111100111111",
    "1110111111110001",
    "1111000011000001",
    "1111000110100101",
    "1111001010010011",
    "1111001110000000",
    "1111010001100010",
    "1111010100101010",
    "1111010111001000",
    "1111011000101000",
    "1111011000111110",
    "1111010111111111",
    "1111010101110001",
    "1111010010100100",
    "1111001110110110",
    "1111001011001110",
    "1111001000010101",
    "1111000110101101",
    "1111000110101101",
    "1111001000010110",
    "1111001011010011",
    "1111001111001010",
    "1111010011010111",
    "1111010111011101",
    "1111011011001010",
    "1111011110011001",
    "1111100001001111",
    "1111100011110110",
    "1111100110011100",
    "1111101001001101",
    "1111101100001111",
    "1111101111100010",
    "1111110011000000",
    "1111110110011000",
    "1111111001011100",
    "1111111011111000",
    "1111111101100010",
    "1111111110010001",
    "1111111101111000",
    "1111111100001101",
    "1111111001001011",
    "1111110100111011",
    "1111101111111011",
    "1111101010111000",
    "1111100110101000",
    "1111100011111000",
    "1111100010111110",
    "1111100011111110",
    "1111100110100000",
    "1111101010000011",
    "1111101101111111",
    "1111110001110101",
    "1111110101001110",
    "1111110111111101",
    "1111111010000110",
    "1111111011110110",
    "1111111101100110",
    "1111111111110001",
    "1111111101001010",
    "1111111000111110",
    "1111110011011010",
    "1111101100011110",
    "1111100100010101",
    "1111011011011001",
    "1111010010010000",
    "1111001001100011",
    "1111000001111000",
    "1110111011110010",
    "1110110111100101",
    "1110110101100100",
    "1110110101110001",
    "1110111000010110",
    "1110111101010010",
    "1111000100011111",
    "1111001101101000",
    "1111011000001011",
    "1111100011001111",
    "1111101101110010",
    "1111110110111010",
    "1111111101111000",
    "1111111101011111",
    "1111111011000111",
    "1111111010011100",
    "1111111010110100",
    "1111111011100110",
    "1111111100010100",
    "1111111100101010",
    "1111111100011101",
    "1111111011101110",
    "1111111010011111",
    "1111111000111010",
    "1111110111001111",
    "1111110101101101",
    "1111110100101001",
    "1111110100010101",
    "1111110101000001",
    "1111110110110111",
    "1111111001111011",
    "1111111110001001",
    "1111111100101000",
    "1111110110110101",
    "1111110000111001",
    "1111101011011000",
    "1111100110110110",
    "1111100011101110",
    "1111100010001101",
    "1111100010001111",
    "1111100011011010",
    "1111100101001101",
    "1111100110111100",
    "1111101000000111",
    "1111101000010001",
    "1111100111010010",
    "1111100101010000",
    "1111100010010100",
    "1111011110101001",
    "1111011010010011",
    "1111010101010010",
    "1111001111100110",
    "1111001001011001",
    "1111000010111110",
    "1110111100101101",
    "1110110111000011",
    "1110110010001111",
    "1110101110010010",
    "1110101010110101",
    "1110100111010011",
    "1110100011010000",
    "1110011110011100",
    "1110011001000100",
    "1110010011101100",
    "1110001111000000",
    "1110001011100110",
    "1110001001101011",
    "1110001001000100",
    "1110001001011110",
    "1110001010110000",
    "1110001100111111",
    "1110010000100001",
    "1110010101110001",
    "1110011100111111",
    "1110100110001000",
    "1110110000100111",
    "1110111011101111",
    "1111000110011011",
    "1111001111110110",
    "1111010111010110",
    "1111011100101110",
    "1111100000001101",
    "1111100010011010",
    "1111100100000000",
    "1111100101100101",
    "1111100111100001",
    "1111101001101111",
    "1111101011111011",
    "1111101101101111",
    "1111101110111001",
    "1111101111010000",
    "1111101110110001",
    "1111101101011011",
    "1111101011000110",
    "1111100111100100",
    "1111100010101100",
    "1111011100010111",
    "1111010100110110",
    "1111001100011011",
    "1111000011100100",
    "1110111010101101",
    "1110110010001010",
    "1110101010001011",
    "1110100010111101",
    "1110011100101000",
    "1110010111010001",
    "1110010010111101",
    "1110001111101011",
    "1110001101100001",
    "1110001100100101",
    "1110001101000010",
    "1110001111000010",
    "1110010010101110",
    "1110011000010101",
    "1110100000000010",
    "1110101010000110",
    "1110110110100101",
    "1111000101010010",
    "1111010101010010",
    "1111100101010011",
    "1111110011111110",
    "1111111111110110",
    "1111110110110101",
    "1111110000110110",
    "1111101101001110",
    "1111101011000000",
    "1111101001010101",
    "1111100111101001",
    "1111100101101100",
    "1111100011011100",
    "1111100000111101",
    "1111011110010001",
    "1111011011011011",
    "1111011000011011",
    "1111010101011011",
    "1111010010101100",
    "1111010000011111",
    "1111001111000101",
    "1111001110100001",
    "1111001110101011",
    "1111001111010111",
    "1111010000010100",
    "1111010001011001",
    "1111010010100001",
    "1111010011100001",
    "1111010100001010",
    "1111010100000110",
    "1111010010111011",
    "1111010000010101",
    "1111001100001100",
    "1111000110100101",
    "1110111111111000",
    "1110111000101101",
    "1110110001110011",
    "1110101011110000",
    "1110100110111001",
    "1110100011010111",
    "1110100001000010",
    "1110011111101001",
    "1110011110111111",
    "1110011110111111",
    "1110011111100100",
    "1110100000110011",
    "1110100010101001",
    "1110100101000000",
    "1110100111101101",
    "1110101010100101",
    "1110101101010111",
    "1110110000000000",
    "1110110010011101",
    "1110110100110100",
    "1110110111011011",
    "1110111010111100",
    "1111000000011110",
    "1111001001001100",
    "1111010110000011",
    "1111100111000101",
    "1111111011001111",
    "1111101111010110",
    "1111011011000111",
    "1111001010001110",
    "1110111101111101",
    "1110110110011010",
    "1110110010100110",
    "1110110001000000",
    "1110110000010111",
    "1110101111111101",
    "1110101111110000",
    "1110110000001101",
    "1110110001101110",
    "1110110100011010",
    "1110110111111010",
    "1110111011100000",
    "1110111110011011",
    "1111000000001100",
    "1111000000101110",
    "1111000000010101",
    "1110111111011001",
    "1110111110001001",
    "1110111100101110",
    "1110111011001110",
    "1110111001100111",
    "1110111000000001",
    "1110110110101111",
    "1110110110010011",
    "1110110111010101",
    "1110111001111101",
    "1110111101111011",
    "1111000010011100",
    "1111000110010011",
    "1111001000100101",
    "1111001000101101",
    "1111000110110010",
    "1111000011011111",
    "1110111111110110",
    "1110111101000000",
    "1110111011110010",
    "1110111100110000",
    "1111000000000111",
    "1111000101110110",
    "1111001101101001",
    "1111010111000011",
    "1111100001011100",
    "1111101100001010",
    "1111110110011110",
    "1111111111101101",
    "1111111000101111",
    "1111110011011001",
    "1111110000010111",
    "1111101111100001",
    "1111110000011100",
    "1111110010100011",
    "1111110101001001",
    "1111110111100011",
    "1111111001010100",
    "1111111010001010",
    "1111111010001110",
    "1111111001101110",
    "1111111000111111",
    "1111111000010000",
    "1111110111101010",
    "1111110111001000",
    "1111110110100011",
    "1111110101101010",
    "1111110100001110",
    "1111110010001010",
    "1111101111100001",
    "1111101100100000",
    "1111101001011111",
    "1111100110111010",
    "1111100101000110",
    "1111100100010101",
    "1111100100100111",
    "1111100101110110",
    "1111100111101010",
    "1111101001101000",
    "1111101011001010",
    "1111101011101000",
    "1111101010011001",
    "1111100111000010",
    "1111100001010101",
    "1111011001011001",
    "1111001111100001",
    "1111000100000101",
    "1110110111100011",
    "1110101010100011",
    "1110011101101000",
    "1110010001011010",
    "1110000110100100",
    "1101111101011011",
    "1101110110001011",
    "1101110000110000",
    "1101101100110111",
    "1101101010001111",
    "1101101000110100",
    "1101101000100101",
    "1101101001101011",
    "1101101100000111",
    "1101101111101001",
    "1101110011111110",
    "1101111000101101",
    "1101111101101000",
    "1110000010101110",
    "1110001000011000",
    "1110001111000101",
    "1110010111010101",
    "1110100001010101",
    "1110101100110111",
    "1110111001010000",
    "1111000101101100",
    "1111010001011001",
    "1111011011100011",
    "1111100011101111",
    "1111101001110001",
    "1111101101110000",
    "1111101111111111",
    "1111110000110111",
    "1111110000110110",
    "1111110000011101",
    "1111110000001100",
    "1111110000010011",
    "1111110000111010",
    "1111110001111111",
    "1111110011011110",
    "1111110101010010",
    "1111110111011100",
    "1111111001111101",
    "1111111100110101",
    "1111111111111100",
    "1111111100111111",
    "1111111010100101",
    "1111111001011001",
    "1111111001111000",
    "1111111100000110",
    "1111111111101000",
    "1111111100010110",
    "1111111000111010",
    "1111110110110111",
    "1111110110100001",
    "1111110111101100",
    "1111111001101010",
    "1111111011100101",
    "1111111100101100",
    "1111111100100001",
    "1111111010111010",
    "1111110111111111",
    "1111110100000100",
    "1111101111100010",
    "1111101010110000",
    "1111100110001001",
    "1111100010001010",
    "1111011111000100",
    "1111011101001010",
    "1111011100100001",
    "1111011101000000",
    "1111011110010001",
    "1111011111110110",
    "1111100001011010",
    "1111100010100111",
    "1111100011011100",
    "1111100011111100",
    "1111100100010111",
    "1111100100110111",
    "1111100101100101",
    "1111100110011101",
    "1111100111011000",
    "1111101000010001",
    "1111101001000001",
    "1111101001101100",
    "1111101010100000",
    "1111101011110000",
    "1111101101110011",
    "1111110000101100",
    "1111110100001101",
    "1111110111110001",
    "1111111010101001",
    "1111111100001100",
    "1111111100001001",
    "1111111010101111",
    "1111111000100111",
    "1111110110100110",
    "1111110101010101",
    "1111110101001000",
    "1111110110000000",
    "1111110111101111",
    "1111111010001111",
    "1111111101011111",
    "1111111110010011",
    "1111111001001001",
    "1111110011000110",
    "1111101100100000",
    "1111100110000000",
    "1111100000010111",
    "1111011100010100",
    "1111011010011101",
    "1111011010111101",
    "1111011101101101",
    "1111100010001011",
    "1111100111101101",
    "1111101101100011",
    "1111110011001000",
    "1111111000001010",
    "1111111100100010",
    "1111111111101110",
    "1111111100110011",
    "1111111010101110",
    "1111111001100010",
    "1111111001000110",
    "1111111001001001",
    "1111111001001111",
    "1111111001000111",
    "1111111000101000",
    "1111110111111101",
    "1111110111011111",
    "1111110111101011",
    "1111111000111011",
    "1111111011010111",
    "1111111110110110",
    "1111111100111001",
    "1111111000011011",
    "1111110100000100",
    "1111110000001011",
    "1111101100111000",
    "1111101010010000",
    "1111101000011101",
    "1111100111101110",
    "1111101000010101",
    "1111101010100010",
    "1111101110010101",
    "1111110011011101",
    "1111111001011000",
    "1111111111010101",
    "1111111011011001",
    "1111110111011000",
    "1111110100110001",
    "1111110011011101",
    "1111110011000110",
    "1111110011010100",
    "1111110011110011",
    "1111110100010111",
    "1111110100111101",
    "1111110101100010",
    "1111110110000010",
    "1111110110011100",
    "1111110110101011",
    "1111110110110111",
    "1111110111001100",
    "1111110111111000",
    "1111111001001110",
    "1111111011010101",
    "1111111110010110",
    "1111111101101100",
    "1111111000110101",
    "1111110010111110",
    "1111101011111100",
    "1111100011100110",
    "1111011001110010",
    "1111001110110000",
    "1111000011001000",
    "1110110111111111",
    "1110101110100001",
    "1110100111110001",
    "1110100100010000",
    "1110100011111000",
    "1110100101111110",
    "1110101001101101",
    "1110101110011001",
    "1110110011101010",
    "1110111001011110",
    "1110111111111000",
    "1111000110110100",
    "1111001101111010",
    "1111010100101001",
    "1111011010011000",
    "1111011110101101",
    "1111100001011111",
    "1111100010111011",
    "1111100011010101",
    "1111100011000101",
    "1111100010011101",
    "1111100001101110",
    "1111100000111101",
    "1111100000001000",
    "1111011111010110",
    "1111011110100001",
    "1111011101101011",
    "1111011100110111",
    "1111011100000111",
    "1111011011011011",
    "1111011010101111",
    "1111011001101111",
    "1111011000000001",
    "1111010101001101",
    "1111010000111110",
    "1111001011010100",
    "1111000100011000",
    "1110111100101000",
    "1110110100100100",
    "1110101100110010",
    "1110100101110010",
    "1110100000000011",
    "1110011011110011",
    "1110011001000110",
    "1110010111110100",
    "1110010111101111",
    "1110011000101101",
    "1110011010100101",
    "1110011101011110",
    "1110100001011010",
    "1110100110011101",
    "1110101100011110",
    "1110110011001111",
    "1110111010011110",
    "1111000001111011",
    "1111001001011001",
    "1111010000101011",
    "1111010111100000",
    "1111011101101000",
    "1111100010101001",
    "1111100110010011",
    "1111101000100010",
    "1111101001100010",
    "1111101001110001",
    "1111101001110010",
    "1111101010001001",
    "1111101011001100",
    "1111101101000010",
    "1111101111100111",
    "1111110010101111",
    "1111110110001101",
    "1111111001110101",
    "1111111101100001",
    "1111111110110011",
    "1111111011001101",
    "1111110111101100",
    "1111110100001110",
    "1111110000101100",
    "1111101101000000",
    "1111101001000010",
    "1111100100101010",
    "1111011111110011",
    "1111011010011110",
    "1111010100110100",
    "1111001111001000",
    "1111001001111001",
    "1111000101100100",
    "1111000010011001",
    "1111000000011100",
    "1110111111010111",
    "1110111110101110",
    "1110111101111011",
    "1110111100101000",
    "1110111010101111",
    "1110111000010110",
    "1110110101111011",
    "1110110011110011",
    "1110110010010010",
    "1110110001100001",
    "1110110001011111",
    "1110110010000010",
    "1110110010111011",
    "1110110100000001",
    "1110110101010000",
    "1110110110100111",
    "1110111000001001",
    "1110111001111101",
    "1110111100000111",
    "1110111110111111",
    "1111000011011010",
    "1111001010110000",
    "1111010110011000",
    "1111100110101111",
    "1111111011001000",
    "1111101110010100",
    "1111011000011101",
    "1111000110001000",
    "1110111001011000",
    "1110110010100100",
    "1110110000100100",
    "1110110001010010",
    "1110110010101001",
    "1110110011010000",
    "1110110010110001",
    "1110110001100010",
    "1110110000010101",
    "1110101111101110",
    "1110101111110000",
    "1110110000000011",
    "1110110000000101",
    "1110101111100001",
    "1110101110010111",
    "1110101100111111",
    "1110101011101111",
    "1110101010110111",
    "1110101010011001",
    "1110101010010011",
    "1110101010011000",
    "1110101010100011",
    "1110101010110010",
    "1110101011001010",
    "1110101011111000",
    "1110101101000010",
    "1110101110101001",
    "1110110000101100",
    "1110110011000101",
    "1110110101101010",
    "1110111000011010",
    "1110111011001010",
    "1110111101111111",
    "1111000000111101",
    "1111000100001110",
    "1111000111111110",
    "1111001100001111",
    "1111010001000111",
    "1111010110011101",
    "1111011100000101",
    "1111100001110000",
    "1111100111000100",
    "1111101011110011",
    "1111101111101101",
    "1111110010101101",
    "1111110100110010",
    "1111110110000001",
    "1111110110101000",
    "1111110110101111",
    "1111110110100000",
    "1111110110000100",
    "1111110101100100",
    "1111110101010001",
    "1111110101100000",
    "1111110110100001",
    "1111111000011010",
    "1111111011001000",
    "1111111110011101",
    "1111111101110111",
    "1111111010001001",
    "1111110110100001",
    "1111110010111010",
    "1111101111000101",
    "1111101010110100",
    "1111100110000001",
    "1111100000110110",
    "1111011011110000",
    "1111010111010101",
    "1111010100000101",
    "1111010010001111",
    "1111010001101001",
    "1111010001110011",
    "1111010010000011",
    "1111010001110000",
    "1111010000100110",
    "1111001110100011",
    "1111001011110000",
    "1111001000011110",
    "1111000100110110",
    "1111000000111011",
    "1110111100101011",
    "1110111000000100",
    "1110110011010101",
    "1110101110101110",
    "1110101010101101",
    "1110100111100101",
    "1110100101100000",
    "1110100100011000",
    "1110100011111000",
    "1110100011011010",
    "1110100010011100",
    "1110100000100100",
    "1110011101110101",
    "1110011010101010",
    "1110010111110101",
    "1110010110001001",
    "1110010110001101",
    "1110011000000001",
    "1110011011010100",
    "1110011111100110",
    "1110100100010111",
    "1110101001011011",
    "1110101110110000",
    "1110110100010011",
    "1110111001111001",
    "1110111111000000",
    "1111000011001010",
    "1111000101111011",
    "1111000111000110",
    "1111000110111001",
    "1111000101101110",
    "1111000100001110",
    "1111000010111110",
    "1111000010010111",
    "1111000010011101",
    "1111000011001010",
    "1111000100001000",
    "1111000101000001",
    "1111000101100101",
    "1111000101101100",
    "1111000101010111",
    "1111000100100111",
    "1111000011011111",
    "1111000010000000",
    "1111000000010010",
    "1110111110011110",
    "1110111100111111",
    "1110111100010001",
    "1110111100110010",
    "1110111110110101",
    "1111000010010111",
    "1111000110111100",
    "1111001011110101",
    "1111010000001101",
    "1111010011011010",
    "1111010101000000",
    "1111010101000001",
    "1111010011101110",
    "1111010001100001",
    "1111001110110110",
    "1111001100000001",
    "1111001001000111",
    "1111000110010110",
    "1111000011110100",
    "1111000001101100",
    "1111000000001010",
    "1110111111011110",
    "1110111111110101",
    "1111000001001101",
    "1111000011100110",
    "1111000110101100",
    "1111001010001110",
    "1111001101111010",
    "1111010001011110",
    "1111010100110111",
    "1111011000000011",
    "1111011010111111",
    "1111011101101011",
    "1111100000001000",
    "1111100010011100",
    "1111100100110011",
    "1111100111100000",
    "1111101010110010",
    "1111101110101100",
    "1111110011000001",
    "1111110111011000",
    "1111111011001111",
    "1111111110000011",
    "1111111111011001",
    "1111111110111101",
    "1111111100100100",
    "1111111000010000",
    "1111110010010011",
    "1111101011010010",
    "1111100100000011",
    "1111011101100110",
    "1111011000110101",
    "1111010110011010",
    "1111010110100000",
    "1111011001000001",
    "1111011101010111",
    "1111100010111001",
    "1111101000111000",
    "1111101110101011",
    "1111110011111100",
    "1111111000100001",
    "1111111100100001",
    "1111111111110000",
    "1111111100000110",
    "1111111000001110",
    "1111110011111110",
    "1111101111010001",
    "1111101010000010",
    "1111100100001110",
    "1111011101110111",
    "1111010111000011",
    "1111010000001100",
    "1111001001101101",
    "1111000100001110",
    "1111000000010010",
    "1110111110010100",
    "1110111110101011",
    "1111000001100001",
    "1111000110110111",
    "1111001110100011",
    "1111010111111111",
    "1111100010011001",
    "1111101100101001",
    "1111110101101010",
    "1111111100100011",
    "1111111110111101",
    "1111111100110101",
    "1111111100011011",
    "1111111100111101",
    "1111111101110000",
    "1111111110010111",
    "1111111110101000",
    "1111111110100101",
    "1111111110010011",
    "1111111101110101",
    "1111111101001010",
    "1111111100001110",
    "1111111011000000",
    "1111111001100101",
    "1111111000001010",
    "1111110110111111",
    "1111110110010100",
    "1111110110010011",
    "1111110110111111",
    "1111111000011000",
    "1111111010010110",
    "1111111100110010",
    "1111111111100001",
    "1111111101100001",
    "1111111010100011",
    "1111110111101001",
    "1111110100111110",
    "1111110010101011",
    "1111110000110110",
    "1111101111100010",
    "1111101110101110",
    "1111101110010001",
    "1111101101111111",
    "1111101101101000",
    "1111101100111110",
    "1111101011110001",
    "1111101001110010",
    "1111100110101111",
    "1111100010011100",
    "1111011100110011",
    "1111010110000000",
    "1111001110010100",
    "1111000110001001",
    "1110111101111010",
    "1110110101110111",
    "1110101110010010",
    "1110100111001011",
    "1110100000011110",
    "1110011010001001",
    "1110010100001101",
    "1110001110111000",
    "1110001010011001",
    "1110000111000110",
    "1110000101010011",
    "1110000101001101",
    "1110000110101000",
    "1110001001010101",
    "1110001100110011",
    "1110010000101100",
    "1110010100110001",
    "1110011001000010",
    "1110011101101000",
    "1110100010110100",
    "1110101000101101",
    "1110101111010001",
    "1110110110010011",
    "1110111101100110",
    "1111000100111011",
    "1111001100000100",
    "1111010010111001",
    "1111011001011011",
    "1111011111100011",
    "1111100101010000",
    "1111101010011010",
    "1111101110110110",
    "1111110010010100",
    "1111110100100110",
    "1111110101100010",
    "1111110101000101",
    "1111110011001101",
    "1111101111111111",
    "1111101011010001",
    "1111100100110110",
    "1111011100011110",
    "1111010010001101",
    "1111000110011010",
    "1110111001111010",
    "1110101101101110",
    "1110100010111001",
    "1110011010000010",
    "1110010011011010",
    "1110001110110001",
    "1110001011101010",
    "1110001001100111",
    "1110001000010011",
    "1110000111101111",
    "1110001000000001",
    "1110001001010101",
    "1110001011110101",
    "1110001111100110",
    "1110010100100010",
    "1110011010100010",
    "1110100001100111",
    "1110101001111001",
    "1110110011100010",
    "1110111110101011",
    "1111001011000001",
    "1111011000000001",
    "1111100100111011",
    "1111110000111101",
    "1111111011100101",
    "1111111011010011",
    "1111110011100100",
    "1111101100110011",
    "1111100110101110",
    "1111100001001111",
    "1111011100100011",
    "1111011000111111",
    "1111010110110110",
    "1111010110001000",
    "1111010110101100",
    "1111011000000110",
    "1111011001110111",
    "1111011011100110",
    "1111011101000101",
    "1111011110001101",
    "1111011110111010",
    "1111011111000000",
    "1111011110011100",
    "1111011101001001",
    "1111011011000110",
    "1111011000100010",
    "1111010101101110",
    "1111010010111001",
    "1111010000010001",
    "1111001101110010",
    "1111001011010100",
    "1111001000101010",
    "1111000101100101",
    "1111000001111001",
    "1110111101100110",
    "1110111000110000",
    "1110110011100111",
    "1110101110100100",
    "1110101010000001",
    "1110100110010101",
    "1110100011101111",
    "1110100010010100",
    "1110100001111000",
    "1110100010010000",
    "1110100011001000",
    "1110100100010010",
    "1110100101100101",
    "1110100111000001",
    "1110101000101000",
    "1110101010100000",
    "1110101100101110",
    "1110101111010111",
    "1110110010011001",
    "1110110101110010",
    "1110111001100000",
    "1110111101100100",
    "1111000010001101",
    "1111000111111110",
    "1111001111101100",
    "1111011010001100",
    "1111100111110101",
    "1111111000010101",
    "1111110101001010",
    "1111100010010010",
    "1111010000110110",
    "1111000010100100",
    "1110111000011010",
    "1110110010100001",
    "1110110000001010",
    "1110110000010001",
    "1110110001101100",
    "1110110011101010",
    "1110110101110010",
    "1110111000000001",
    "1110111010011101",
    "1110111100111100",
    "1110111111001100",
    "1111000000101100",
    "1111000001001100",
    "1111000000011111",
    "1110111110110101",
    "1110111100100001",
    "1110111001111010",
    "1110110111010001",
    "1110110100101110",
    "1110110010010010",
    "1110101111111011",
    "1110101101101110",
    "1110101011110010",
    "1110101010010110",
    "1110101001101010",
    "1110101001110101",
    "1110101010111100",
    "1110101101000000",
    "1110110000000000",
    "1110110011111110",
    "1110111000110100",
    "1110111110011100",
    "1111000100101001",
    "1111001011000111",
    "1111010001100001",
    "1111010111100010",
    "1111011100110010",
    "1111100000111110",
    "1111100100000011",
    "1111100110000001",
    "1111100111010001",
    "1111101000010001",
    "1111101001100010",
    "1111101011011110",
    "1111101110001101",
    "1111110001100111",
    "1111110101010111",
    "1111111001001000",
    "1111111100101010",
    "1111111111111100",
    "1111111100111110",
    "1111111010000000",
    "1111110111000100",
    "1111110100001101",
    "1111110001101100",
    "1111101111110100",
    "1111101110110011",
    "1111101110101110",
    "1111101111011000",
    "1111110000011001",
    "1111110001010011",
    "1111110001101110",
    "1111110001011110",
    "1111110000100110",
    "1111101111011001",
    "1111101110001100",
    "1111101101010000",
    "1111101100101011",
    "1111101100100000",
    "1111101100100111",
    "1111101100110101",
    "1111101100111111",
    "1111101100110101",
    "1111101100000111",
    "1111101010011101",
    "1111100111100010",
    "1111100010111110",
    "1111011100100101",
    "1111010100001011",
    "1111001001111001",
    "1110111101111010",
    "1110110000110011",
    "1110100011010011",
    "1110010110010110",
    "1110001010110100",
    "1110000001010100",
    "1101111010000100",
    "1101110101000001",
    "1101110001110001",
    "1101101111111101",
    "1101101111001111",
    "1101101111011010",
    "1101110000011110",
    "1101110010010000",
    "1101110100101100",
    "1101110111100101",
    "1101111010110111",
    "1101111110100011",
    "1110000010110011",
    "1110000111110010",
    "1110001101101101",
    "1110010100100100",
    "1110011100010011",
    "1110100100100100",
    "1110101101000000",
    "1110110101010000",
    "1110111100111010",
    "1111000011101110",
    "1111001001100011",
    "1111001110011100",
    "1111010010100001",
    "1111010110000100",
    "1111011001011000",
    "1111011100101000",
    "1111100000000011",
    "1111100011101110",
    "1111100111100110",
    "1111101011100011",
    "1111101111011000",
    "1111110010111110",
    "1111110110001101",
    "1111111001001000",
    "1111111011110000",
    "1111111110001011",
    "1111111111100110",
    "1111111101110000",
    "1111111100100001",
    "1111111100001101",
    "1111111101000001",
    "1111111110111010",
    "1111111110011100",
    "1111111011101110",
    "1111111001101000",
    "1111111000101011",
    "1111111001000101",
    "1111111010100111",
    "1111111100101010",
    "1111111110011111",
    "1111111111011010",
    "1111111110111010",
    "1111111100101110",
    "1111111000111000",
    "1111110011101001",
    "1111101101100101",
    "1111100111010111",
    "1111100001101100",
    "1111011101001110",
    "1111011010010110",
    "1111011001010001",
    "1111011001111101",
    "1111011100001110",
    "1111011111101001",
    "1111100011110110",
    "1111101000010100",
    "1111101100100011",
    "1111110000000100",
    "1111110010100001",
    "1111110011100111",
    "1111110011010100",
    "1111110001101001",
    "1111101110110011",
    "1111101011001010",
    "1111100111001000",
    "1111100011001111",
    "1111100000000000",
    "1111011101110111",
    "1111011101001010",
    "1111011101111111",
    "1111100000001100",
    "1111100011011101",
    "1111100111001111",
    "1111101010111110",
    "1111101110001011",
    "1111110000100011",
    "1111110010000110",
    "1111110011000001",
    "1111110011110000",
    "1111110100101100",
    "1111110110001010",
    "1111111000010001",
    "1111111011000100",
    "1111111110100100",
    "1111111101001001",
    "1111111000000010",
    "1111110010000110",
    "1111101011100100",
    "1111100100111001",
    "1111011110110001",
    "1111011001111001",
    "1111010110110001",
    "1111010101101110",
    "1111010110111001",
    "1111011010001110",
    "1111011111100100",
    "1111100110101101",
    "1111101111001110",
    "1111111000100111",
    "1111111101110110",
    "1111110101001100",
    "1111101110010010",
    "1111101001110100",
    "1111101000000111",
    "1111101000111110",
    "1111101011101111",
    "1111101111100001",
    "1111110011011001",
    "1111110110110001",
    "1111111001011001",
    "1111111011011101",
    "1111111101010010",
    "1111111111010110",
    "1111111110000101",
    "1111111011000001",
    "1111110111101101",
    "1111110100100010",
    "1111110001111101",
    "1111110000010001",
    "1111101111100010",
    "1111101111101011",
    "1111110000011100",
    "1111110001100100",
    "1111110010111001",
    "1111110100011001",
    "1111110110000111",
    "1111111000000110",
    "1111111010011000",
    "1111111100111001",
    "1111111111011101",
    "1111111110000110",
    "1111111100000001",
    "1111111010010011",
    "1111111000110011",
    "1111110111001111",
    "1111110101011010",
    "1111110011001010",
    "1111110000101001",
    "1111101110000111",
    "1111101011111010",
    "1111101010011010",
    "1111101001110100",
    "1111101010001010",
    "1111101011011010",
    "1111101101100000",
    "1111110000011000",
    "1111110100000110",
    "1111111000101101",
    "1111111110001100",
    "1111111011100011",
    "1111110100110110",
    "1111101101111010",
    "1111100110111011",
    "1111011111111011",
    "1111011000111001",
    "1111010001110000",
    "1111001010100010",
    "1111000011011100",
    "1110111100110011",
    "1110110111000100",
    "1110110010101011",
    "1110110000000000",
    "1110101111001111",
    "1110110000001010",
    "1110110010010101",
    "1110110101001000",
    "1110111000001011",
    "1110111011011000",
    "1110111111000000",
    "1111000011100001",
    "1111001001001100",
    "1111001111111011",
    "1111010111001000",
    "1111011101111111",
    "1111100011110100",
    "1111101000001111",
    "1111101011001001",
    "1111101100110011",
    "1111101101011011",
    "1111101101001111",
    "1111101100010100",
    "1111101010101010",
    "1111101000001110",
    "1111100101000000",
    "1111100001000011",
    "1111011100100000",
    "1111010111100000",
    "1111010010010100",
    "1111001101000010",
    "1111000111101101",
    "1111000010010100",
    "1110111100101010",
    "1110110110101111",
    "1110110000100111",
    "1110101010100101",
    "1110100101000001",
    "1110100000001111",
    "1110011100011001",
    "1110011001011011",
    "1110010111000001",
    "1110010100110111",
    "1110010010110100",
    "1110010000111110",
    "1110001111110000",
    "1110001111101011",
    "1110010001001101",
    "1110010100101010",
    "1110011010001001",
    "1110100001101011",
    "1110101010111111",
    "1110110101110110",
    "1111000001101110",
    "1111001101111011",
    "1111011001101010",
    "1111100100000101",
    "1111101100100000",
    "1111110010100000",
    "1111110101111000",
    "1111110110110001",
    "1111110101100011",
    "1111110010101100",
    "1111101110110101",
    "1111101010101100",
    "1111100110111111",
    "1111100100011010",
    "1111100011011100",
    "1111100100010010",
    "1111100110111000",
    "1111101010111001",
    "1111101111110100",
    "1111110101000010",
    "1111111010000101",
    "1111111110101100",
    "1111111101000100",
    "1111111001000010",
    "1111110100110110",
    "1111110000010101",
    "1111101011011100",
    "1111100110010010",
    "1111100001000011",
    "1111011011111100",
    "1111010110111111",
    "1111010010010100",
    "1111001101111101",
    "1111001010001011",
    "1111000111001001",
    "1111000100111110",
    "1111000011011100",
    "1111000010001011",
    "1111000000110000",
    "1110111110101011",
    "1110111011110111",
    "1110111000011110",
    "1110110101000011",
    "1110110010000110",
    "1110110000001100",
    "1110101111011110",
    "1110101111111011",
    "1110110001010010",
    "1110110011001010",
    "1110110101010000",
    "1110110111011010",
    "1110111001100000",
    "1110111011100101",
    "1110111101101011",
    "1110111111111010",
    "1111000010011001",
    "1111000101101010",
    "1111001010110101",
    "1111010011001011",
    "1111011111101000",
    "1111110000001011",
    "1111111100010011",
    "1111100111111001",
    "1111010101001011",
    "1111000110011000",
    "1110111100101101",
    "1110110111111110",
    "1110110110110010",
    "1110110111010001",
    "1110110111110001",
    "1110110111010011",
    "1110110101110001",
    "1110110011101110",
    "1110110001111001",
    "1110110000110101",
    "1110110000100001",
    "1110110000101011",
    "1110110000110101",
    "1110110000100110",
    "1110101111111010",
    "1110101110110011",
    "1110101101011110",
    "1110101011111101",
    "1110101010010001",
    "1110101000011011",
    "1110100110100000",
    "1110100100100111",
    "1110100010111001",
    "1110100001101011",
    "1110100001001111",
    "1110100001111011",
    "1110100011110100",
    "1110100110111110",
    "1110101011010001",
    "1110110000100111",
    "1110110110110111",
    "1110111101110000",
    "1111000100111011",
    "1111001011110011",
    "1111010001110011",
    "1111010110011111",
    "1111011001101011",
    "1111011011100110",
    "1111011100101110",
    "1111011101101001",
    "1111011110110110",
    "1111100000100011",
    "1111100010101100",
    "1111100101000101",
    "1111100111011111",
    "1111101001101101",
    "1111101011100110",
    "1111101101000111",
    "1111101110010000",
    "1111101110111111",
    "1111101111011110",
    "1111101111111010",
    "1111110000101111",
    "1111110010011001",
    "1111110101010001",
    "1111111001010111",
    "1111111110011100",
    "1111111011111100",
    "1111110110011101",
    "1111110001011101",
    "1111101101001001",
    "1111101001100011",
    "1111100110100101",
    "1111100100001010",
    "1111100010010000",
    "1111100000111000",
    "1111100000000000",
    "1111011111011100",
    "1111011110111000",
    "1111011101111010",
    "1111011100001100",
    "1111011001100011",
    "1111010110000011",
    "1111010010000000",
    "1111001101110010",
    "1111001001101010",
    "1111000101110010",
    "1111000010000011",
    "1110111110001100",
    "1110111001111101",
    "1110110101010101",
    "1110110000011111",
    "1110101011101011",
    "1110100111010101",
    "1110100011101100",
    "1110100000111001",
    "1110011110111010",
    "1110011101100100",
    "1110011100100101",
    "1110011011101101",
    "1110011010111010",
    "1110011010010011",
    "1110011010001111",
    "1110011011001001",
    "1110011101010110",
    "1110100000110110",
    "1110100101011010",
    "1110101010011101",
    "1110101111010111",
    "1110110011101001",
    "1110110111000001",
    "1110111001100000",
    "1110111011010001",
    "1110111100100001",
    "1110111101011100",
    "1110111110001010",
    "1110111110101000",
    "1110111110110000",
    "1110111110100001",
    "1110111101111000",
    "1110111101000100",
    "1110111100010011",
    "1110111011111010",
    "1110111100001100",
    "1110111101001110",
    "1110111110111010",
    "1111000001000000",
    "1111000011000110",
    "1111000100110100",
    "1111000101110100",
    "1111000101110110",
    "1111000100111001",
    "1111000011000011",
    "1111000000101110",
    "1110111110011100",
    "1110111100110111",
    "1110111100101011",
    "1110111110010110",
    "1111000001111110",
    "1111000111001011",
    "1111001101000101",
    "1111010010101111",
    "1111010111001001",
    "1111011001101000",
    "1111011001111100",
    "1111011000001100",
    "1111010100110001",
    "1111010000000101",
    "1111001010100101",
    "1111000100101001",
    "1110111110101001",
    "1110111001000110",
    "1110110100100000",
    "1110110001010111",
    "1110110000000010",
    "1110110000101001",
    "1110110011000101",
    "1110110111000110",
    "1110111100010110",
    "1111000010011010",
    "1111001000111111",
    "1111001111110001",
    "1111010110011101",
    "1111011100101101",
    "1111100010010000",
    "1111100110111000",
    "1111101010011000",
    "1111101100101101",
    "1111101101111100",
    "1111101110010100",
    "1111101110010001",
    "1111101110010011",
    "1111101110110101",
    "1111110000000000",
    "1111110001100100",
    "1111110011000001",
    "1111110011110011",
    "1111110011011010",
    "1111110001100111",
    "1111101110011001",
    "1111101001111111",
    "1111100100110110",
    "1111011111100110",
    "1111011010111100",
    "1111010111100000",
    "1111010101101110",
    "1111010101101110",
    "1111010111010110",
    "1111011010001110",
    "1111011101111111",
    "1111100010011101",
    "1111100111100011",
    "1111101101010100",
    "1111110011101100",
    "1111111010011111",
    "1111111110100001",
    "1111110111101000",
    "1111110001000001",
    "1111101010110011",
    "1111100101001000",
    "1111100000001000",
    "1111011011111111",
    "1111011000110101",
    "1111010110101010",
    "1111010101011000",
    "1111010100101010",
    "1111010100010101",
    "1111010100010111",
    "1111010100111100",
    "1111010110011011",
    "1111011001000100",
    "1111011100111000",
    "1111100001101011",
    "1111100110111010",
    "1111101011111100",
    "1111110000010000",
    "1111110011100001",
    "1111110101110000",
    "1111110111001101",
    "1111111000010001",
    "1111111001011000",
    "1111111010110101",
    "1111111100101101",
    "1111111110111010",
    "1111111110110100",
    "1111111100110110",
    "1111111011010101",
    "1111111010010001",
    "1111111001100010",
    "1111111000111110",
    "1111111000011011",
    "1111110111111001",
    "1111110111100001",
    "1111110111011101",
    "1111110111111001",
    "1111111000111001",
    "1111111010010101",
    "1111111011111110",
    "1111111101100001",
    "1111111110101101",
    "1111111111010110",
    "1111111111011010",
    "1111111110111101",
    "1111111110001101",
    "1111111101011101",
    "1111111101000000",
    "1111111101001000",
    "1111111101111111",
    "1111111111101001",
    "1111111101110101",
    "1111111010100111",
    "1111110110110010",
    "1111110010100100",
    "1111101110001100",
    "1111101001110110",
    "1111100101100101",
    "1111100001010100",
    "1111011100111000",
    "1111011000001011",
    "1111010011000011",
    "1111001101100001",
    "1111000111101000",
    "1111000001011010",
    "1110111010111100",
    "1110110100001101",
    "1110101101001111",
    "1110100110000011",
    "1110011110101110",
    "1110010111011010",
    "1110010000010101",
    "1110001001110111",
    "1110000100010011",
    "1101111111111101",
    "1101111101000000",
    "1101111011100011",
    "1101111011101011",
    "1101111101100110",
    "1110000001100010",
    "1110000111101010",
    "1110001111111111",
    "1110011010001110",
    "1110100101110001",
    "1110110001110100",
    "1110111101100011",
    "1111001000010011",
    "1111010001100110",
    "1111011001001100",
    "1111011111000010",
    "1111100011001011",
    "1111100101110111",
    "1111100111011101",
    "1111101000010111",
    "1111101000111110",
    "1111101001100011",
    "1111101010001100",
    "1111101010110001",
    "1111101011000001",
    "1111101010101001",
    "1111101001001111",
    "1111100110011000",
    "1111100001100001",
    "1111011010000111",
    "1111001111111111",
    "1111000011011101",
    "1110110101011111",
    "1110100111011101",
    "1110011010101011",
    "1110010000001100",
    "1110001000010110",
    "1110000010111110",
    "1101111111100110",
    "1101111101101011",
    "1101111100110111",
    "1101111101000101",
    "1101111110100011",
    "1110000001010111",
    "1110000101101001",
    "1110001011010100",
    "1110010010010100",
    "1110011010011000",
    "1110100011010101",
    "1110101101000100",
    "1110110111011111",
    "1111000010011001",
    "1111001101100100",
    "1111011000101000",
    "1111100011001101",
    "1111101101000111",
    "1111110110010000",
    "1111111110101100",
    "1111111001011111",
    "1111110010011100",
    "1111101100010110",
    "1111100111100000",
    "1111100100001011",
    "1111100010011100",
    "1111100010001000",
    "1111100010111001",
    "1111100100001011",
    "1111100101011010",
    "1111100110010000",
    "1111100110011011",
    "1111100101110111",
    "1111100100101110",
    "1111100011000011",
    "1111100001000011",
    "1111011110110101",
    "1111011100100011",
    "1111011010011011",
    "1111011000101000",
    "1111010111010000",
    "1111010110001110",
    "1111010101011000",
    "1111010100011010",
    "1111010010111011",
    "1111010000100100",
    "1111001101001010",
    "1111001000101101",
    "1111000011010101",
    "1110111101010110",
    "1110110111000100",
    "1110110000110110",
    "1110101011000111",
    "1110100110010000",
    "1110100010100111",
    "1110100000011100",
    "1110011111110000",
    "1110100000010100",
    "1110100001110100",
    "1110100011110001",
    "1110100101110100",
    "1110100111101111",
    "1110101001100011",
    "1110101011011001",
    "1110101101011110",
    "1110101111111111",
    "1110110010111110",
    "1110110110010110",
    "1110111010000100",
    "1110111101111111",
    "1111000010001000",
    "1111000110111100",
    "1111001101000111",
    "1111010101010111",
    "1111100000000101",
    "1111101101000011",
    "1111111011010011",
    "1111110110100000",
    "1111101001110000",
    "1111011111010111",
    "1111010111101100",
    "1111010010011100",
    "1111001110111011",
    "1111001100010110",
    "1111001001111111",
    "1111000111011101",
    "1111000100100111",
    "1111000001100010",
    "1110111110011111",
    "1110111011110000",
    "1110111001100101",
    "1110111000001011",
    "1110110111011011",
    "1110110111001101",
    "1110110111010000",
    "1110110111010000",
    "1110110110111100",
    "1110110110001011",
    "1110110100111011",
    "1110110011010011",
    "1110110001100001",
    "1110101111101000",
    "1110101101110000",
    "1110101011111101",
    "1110101010011001",
    "1110101001010000",
    "1110101000110100",
    "1110101001011110",
    "1110101011100000",
    "1110101111000000",
    "1110110011110110",
    "1110111001100101",
    "1110111111101011",
    "1111000101011011",
    "1111001010011011",
    "1111001110011001",
    "1111010001010101",
    "1111010011011101",
    "1111010101000011",
    "1111010110011000",
    "1111010111101101",
    "1111011001010101",
    "1111011011011001",
    "1111011110001001",
    "1111100001110000",
    "1111100110001101",
    "1111101011010101",
    "1111110000111010",
    "1111110110101001",
    "1111111100010011",
    "1111111110010001",
    "1111111001001111",
    "1111110100101101",
    "1111110000111100",
    "1111101110001100",
    "1111101100101111",
    "1111101100100110",
    "1111101101100110",
    "1111101111011010",
    "1111110001101000",
    "1111110011111000",
    "1111110101111011",
    "1111110111100101",
    "1111111000101110",
    "1111111001010010",
    "1111111001001111",
    "1111111000101011",
    "1111110111101100",
    "1111110110011000",
    "1111110100110101",
    "1111110011000111",
    "1111110001001110",
    "1111101111001011",
    "1111101100110110",
    "1111101010000100",
    "1111100110011110",
    "1111100001101100",
    "1111011011010110",
    "1111010011010010",
    "1111001001101010",
    "1110111110110110",
    "1110110011100010",
    "1110101000011010",
    "1110011110000111",
    "1110010101010000",
    "1110001110001100",
    "1110001001000001",
    "1110000101101010",
    "1110000011110011",
    "1110000010111011",
    "1110000010100100",
    "1110000010010100",
    "1110000001111101",
    "1110000001011110",
    "1110000000111001",
    "1110000000010111",
    "1101111111111111",
    "1101111111111011",
    "1110000000011010",
    "1110000001111000",
    "1110000100100111",
    "1110001000111010",
    "1110001110110000",
    "1110010101110100",
    "1110011101100110",
    "1110100101100010",
    "1110101101010010",
    "1110110100100100",
    "1110111011001111",
    "1111000001001101",
    "1111000110011000",
    "1111001010101011",
    "1111001110001111",
    "1111010001001111",
    "1111010100000001",
    "1111010111000011",
    "1111011010100011",
    "1111011110101101",
    "1111100011010111",
    "1111101000010010",
    "1111101101001100",
    "1111110001111001",
    "1111110110010000",
    "1111111010010001",
    "1111111101111010",
    "1111111110110110",
    "1111111100001111",
    "1111111010011100",
    "1111111001101110",
    "1111111010010010",
    "1111111100001011",
    "1111111111001101",
    "1111111100111101",
    "1111111001000011",
    "1111110101101010",
    "1111110011001110",
    "1111110001111100",
    "1111110001101110",
    "1111110010001010",
    "1111110010110010",
    "1111110011001000",
    "1111110010110111",
    "1111110001111100",
    "1111110000100011",
    "1111101110111100",
    "1111101101011010",
    "1111101100001011",
    "1111101011010001",
    "1111101010101110",
    "1111101010100011",
    "1111101010110000",
    "1111101011011011",
    "1111101100100010",
    "1111101101111110",
    "1111101111011000",
    "1111110000011011",
    "1111110000110010",
    "1111110000010111",
    "1111101111001011",
    "1111101101011010",
    "1111101011010000",
    "1111101000110101",
    "1111100110001001",
    "1111100011010000",
    "1111100000001010",
    "1111011101000100",
    "1111011010001111",
    "1111011000001001",
    "1111010111001000",
    "1111010111011010",
    "1111011000111100",
    "1111011011100110",
    "1111011111000010",
    "1111100010111101",
    "1111100111001011",
    "1111101011101000",
    "1111110000011101",
    "1111110101101111",
    "1111111011100100",
    "1111111110001010",
    "1111110111110010",
    "1111110001100011",
    "1111101011110010",
    "1111100110101100",
    "1111100010011101",
    "1111011111010010",
    "1111011101010110",
    "1111011100110101",
    "1111011101110000",
    "1111011111111011",
    "1111100011000101",
    "1111100110111000",
    "1111101011001011",
    "1111101111111111",
    "1111110101010111",
    "1111111011010010",
    "1111111110011001",
    "1111111000001000",
    "1111110010011010",
    "1111101101110101",
    "1111101010101101",
    "1111101001001111",
    "1111101001010010",
    "1111101010100001",
    "1111101100100000",
    "1111101110110111",
    "1111110001011000",
    "1111110100000110",
    "1111110111001010",
    "1111111010110010",
    "1111111111000101",
    "1111111011111110",
    "1111110110110010",
    "1111110001110011",
    "1111101101100101",
    "1111101010100111",
    "1111101001001100",
    "1111101001010110",
    "1111101010111010",
    "1111101101100100",
    "1111110000111111",
    "1111110100110100",
    "1111111000110000",
    "1111111100100111",
    "1111111111110110",
    "1111111100111001",
    "1111111010100101",
    "1111111000111110",
    "1111110111111000",
    "1111110111000111",
    "1111110110011000",
    "1111110101011011",
    "1111110100001000",
    "1111110010011110",
    "1111110000100011",
    "1111101110011010",
    "1111101100001000",
    "1111101001101101",
    "1111100111001000",
    "1111100100011010",
    "1111100001101110",
    "1111011111010100",
    "1111011101100100",
    "1111011100111010",
    "1111011101101110",
    "1111100000010100",
    "1111100100110011",
    "1111101011001111",
    "1111110011100001",
    "1111111101011100",
    "1111110111001100",
    "1111101010100101",
    "1111011100110010",
    "1111001101111011",
    "1110111110101001",
    "1110101111110011",
    "1110100010100010",
    "1110011000000100",
    "1110010001010000",
    "1110001110011100",
    "1110001111010010",
    "1110010010111101",
    "1110011000010110",
    "1110011110101110",
    "1110100101111011",
    "1110101110000100",
    "1110110111100000",
    "1111000010010111",
    "1111001110001010",
    "1111011001111111",
    "1111100100101100",
    "1111101101010000",
    "1111110011001001",
    "1111110110011111",
    "1111110111111100",
    "1111111000010010",
    "1111111000001100",
    "1111111000000001",
    "1111110111110101",
    "1111110111010111",
    "1111110110001110",
    "1111110011111100",
    "1111110000000110",
    "1111101010011001",
    "1111100010101110",
    "1111011000111111",
    "1111001101011001",
    "1111000000001111",
    "1110110010010101",
    "1110100100101001",
    "1110011000010011",
    "1110001110001001",
    "1110000110101000",
    "1110000001101110",
    "1101111110110101",
    "1101111101010100",
    "1101111100100011",
    "1101111100010011",
    "1101111100110000",
    "1101111110010110",
    "1110000001100001",
    "1110000110101101",
    "1110001110000111",
    "1110010111110101",
    "1110100011111000",
    "1110110010001000",
    "1111000010000110",
    "1111010010110110",
    "1111100011000000",
    "1111110001000011",
    "1111111011110000",
    "1111111101100101",
    "1111111010111010",
    "1111111011011100",
    "1111111110000101",
    "1111111110000111",
    "1111111001110100",
    "1111110101010000",
    "1111110000010011",
    "1111101010111010",
    "1111100101001001",
    "1111011111011010",
    "1111011010010100",
    "1111010110011011",
    "1111010100000110",
    "1111010011011100",
    "1111010100010010",
    "1111010110011000",
    "1111011001101111",
    "1111011110011100",
    "1111100100101100",
    "1111101100100101",
    "1111110101110011",
    "1111111111101001",
    "1111110110101111",
    "1111101110010101",
    "1111100111101110",
    "1111100010111110",
    "1111011111101001",
    "1111011100111111",
    "1111011010001100",
    "1111010110100111",
    "1111010010000011",
    "1111001100101000",
    "1111000110101101",
    "1111000000110001",
    "1110111011001001",
    "1110110110000011",
    "1110110001101100",
    "1110101110001001",
    "1110101011011110",
    "1110101001110000",
    "1110101000111111",
    "1110101001001001",
    "1110101010000100",
    "1110101011100101",
    "1110101101011100",
    "1110101111100001",
    "1110110001110000",
    "1110110100001011",
    "1110110110111110",
    "1110111010001100",
    "1110111101111101",
    "1111000010000110",
    "1111000110011011",
    "1111001010101011",
    "1111001110101011",
    "1111010010100100",
    "1111010110110111",
    "1111011100001110",
    "1111100011010000",
    "1111101100010010",
    "1111110111000001",
    "1111111101001010",
    "1111110001001101",
    "1111100101111110",
    "1111011100000111",
    "1111010011111000",
    "1111001101001100",
    "1111000111101101",
    "1111000011000001",
    "1110111110110101",
    "1110111010111101",
    "1110110111100000",
    "1110110100101001",
    "1110110010100100",
    "1110110001001111",
    "1110110000010111",
    "1110101111100100",
    "1110101110010110",
    "1110101100010111",
    "1110101001100011",
    "1110100110000001",
    "1110100010000101",
    "1110011110001111",
    "1110011011000100",
    "1110011001010101",
    "1110011010000010",
    "1110011110001010",
    "1110100110000110",
    "1110110001011010",
    "1110111110101011",
    "1111001011101000",
    "1111010101111011",
    "1111011011110000",
    "1111011100100110",
    "1111011001001100",
    "1111010011000101",
    "1111001011111101",
    "1111000101010000",
    "1110111111110001",
    "1110111011110011",
    "1110111001011001",
    "1110111000100000",
    "1110111001000110",
    "1110111011000010",
    "1110111110000000",
    "1111000001011110",
    "1111000100110110",
    "1111000111101100",
    "1111001001110100",
    "1111001011011101",
    "1111001101010110",
    "1111010000100110",
    "1111010110011010",
    "1111011111100100",
    "1111101100010010",
    "1111111011110011",
    "1111110011001100",
    "1111100010100010",
    "1111010100000101",
    "1111001001010001",
    "1111000011000000",
    "1111000001010111",
    "1111000011110100",
    "1111001001011011",
    "1111010001000101",
    "1111011001110100",
    "1111100010110011",
    "1111101011010111",
    "1111110010111100",
    "1111111000111111",
    "1111111101000101",
    "1111111110111100",
    "1111111110100110",
    "1111111100010111",
    "1111111000101111",
    "1111110100010100",
    "1111101111100100",
    "1111101010110110",
    "1111100110001110",
    "1111100001100001",
    "1111011100011110",
    "1111010110111001",
    "1111010000101110",
    "1111001010000110",
    "1111000011010111",
    "1110111100111000",
    "1110110110110110",
    "1110110001001111",
    "1110101011110011",
    "1110100110010000",
    "1110100000010111",
    "1110011010001001",
    "1110010011110110",
    "1110001101111111",
    "1110001001010101",
    "1110000110110100",
    "1110000111010001",
    "1110001011000100",
    "1110010010000000",
    "1110011011010110",
    "1110100110000100",
    "1110110001000111",
    "1110111011100011",
    "1111000100110011",
    "1111001100011100",
    "1111010010001111",
    "1111010101111100",
    "1111010111101000",
    "1111010111100101",
    "1111010110010101",
    "1111010100100101",
    "1111010011000101",
    "1111010010001111",
    "1111010010001101",
    "1111010010110001",
    "1111010011011111",
    "1111010011111001",
    "1111010011100001",
    "1111010010000101",
    "1111001111010110",
    "1111001011001100",
    "1111000101100100",
    "1110111110101001",
    "1110110110110100",
    "1110101110110101",
    "1110100111100111",
    "1110100010000110",
    "1110011111000100",
    "1110011110101110",
    "1110100000111011",
    "1110100101010000",
    "1110101011000100",
    "1110110001111000",
    "1110111001010001",
    "1111000001000011",
    "1111001001000111",
    "1111010001010000",
    "1111011001001100",
    "1111100000100011",
    "1111100110111000",
    "1111101011110011",
    "1111101111001011",
    "1111110000111100",
    "1111110001001100",
    "1111110000000001",
    "1111101101011011",
    "1111101001011010",
    "1111100100000001",
    "1111011101100011",
    "1111010110100100",
    "1111001111101100",
    "1111001001110100",
    "1111000101011011",
    "1111000010111101",
    "1111000010010010",
    "1111000011001010",
    "1111000101000110",
    "1111000111101000",
    "1111001010011101",
    "1111001101010110",
    "1111010000001111",
    "1111010011010000",
    "1111010110100010",
    "1111011010001111",
    "1111011110011100",
    "1111100010111110",
    "1111100111011111",
    "1111101011100011",
    "1111101110110001",
    "1111110000111100",
    "1111110010001101",
    "1111110010111001",
    "1111110011100100",
    "1111110100101110",
    "1111110110110011",
    "1111111001110111",
    "1111111101101001",
    "1111111110011010",
    "1111111011001001",
    "1111111001000110",
    "1111111000101000",
    "1111111001101000",
    "1111111011110000",
    "1111111110100011",
    "1111111110010010",
    "1111111011000100",
    "1111110111111001",
    "1111110100111010",
    "1111110010011001",
    "1111110000101110",
    "1111110000001001",
    "1111110000101110",
    "1111110010000110",
    "1111110011111011",
    "1111110101110111",
    "1111110111111000",
    "1111111010000110",
    "1111111100101000",
    "1111111111011110",
    "1111111101100101",
    "1111111010111111",
    "1111111001000000",
    "1111110111101101",
    "1111110110110010",
    "1111110101101010",
    "1111110011101010",
    "1111110000011000",
    "1111101011101111",
    "1111100110000011",
    "1111100000000101",
    "1111011010110000",
    "1111010110111111",
    "1111010101100000",
    "1111010110100000",
    "1111011001100111",
    "1111011110000000",
    "1111100010110001",
    "1111100111001010",
    "1111101010110010",
    "1111101101101000",
    "1111110000000010",
    "1111110010010111",
    "1111110100111101",
    "1111110111111101",
    "1111111011010011",
    "1111111110110010",
    "1111111101110101",
    "1111111010110111",
    "1111111000011101",
    "1111110110101111",
    "1111110101101000",
    "1111110101000011",
    "1111110100110001",
    "1111110100101011",
    "1111110100110100",
    "1111110101010101",
    "1111110110100001",
    "1111111000101010",
    "1111111011111000",
    "1111111111111001",
    "1111111011000011",
    "1111110110000001",
    "1111110001001110",
    "1111101101000011",
    "1111101001101001",
    "1111100111000110",
    "1111100101011000",
    "1111100100011000",
    "1111100011111000",
    "1111100011100111",
    "1111100011010000",
    "1111100010100111",
    "1111100001100010",
    "1111100000001100",
    "1111011110110101",
    "1111011101111000",
    "1111011101101000",
    "1111011110000111",
    "1111011111000000",
    "1111011111110001",
    "1111011111101001",
    "1111011101111111",
    "1111011010010100",
    "1111010100100010",
    "1111001100101010",
    "1111000011001010",
    "1110111000110100",
    "1110101110101101",
    "1110100110000011",
    "1110011111110101",
    "1110011100101101",
    "1110011100110011",
    "1110011111111011",
    "1110100101100101",
    "1110101101001110",
    "1110110110010110",
    "1111000000100100",
    "1111001011010001",
    "1111010101101110",
    "1111011111000000",
    "1111100110010011",
    "1111101011000101",
    "1111101101010001",
    "1111101101010000",
    "1111101011101010",
    "1111101001001111",
    "1111100110100010",
    "1111100011101110",
    "1111100000110000",
    "1111011101010110",
    "1111011001001110",
    "1111010100001011",
    "1111001101111011",
    "1111000110010011",
    "1110111101010001",
    "1110110011001011",
    "1110101000101100",
    "1110011110101101",
    "1110010101111100",
    "1110001110111010",
    "1110001001100011",
    "1110000101100100",
    "1110000010010101",
    "1101111111011010",
    "1101111100101011",
    "1101111010010011",
    "1101111000101000",
    "1101111000000001",
    "1101111000100111",
    "1101111010011000",
    "1101111101010001",
    "1110000001011001",
    "1110000111010101",
    "1110010000001000",
    "1110011100111101",
    "1110101110010100",
    "1111000011011101",
    "1111011010100010",
    "1111110000111000",
    "1111111100000011",
    "1111101110001011",
    "1111100101111100",
    "1111100010101100",
    "1111100010110100",
    "1111100100100100",
    "1111100110100010",
    "1111100111111101",
    "1111101000100110",
    "1111101000101100",
    "1111101000100101",
    "1111101000100111",
    "1111101001000100",
    "1111101010001001",
    "1111101100000010",
    "1111101110111100",
    "1111110010111110",
    "1111110111111011",
    "1111111101010001",
    "1111111101101111",
    "1111111001111110",
    "1111111000000101",
    "1111111000011011",
    "1111111011001001",
    "1111111111111101",
    "1111111001011101",
    "1111110010000010",
    "1111101010011111",
    "1111100011011111",
    "1111011101100001",
    "1111011000101010",
    "1111010100100100",
    "1111010000101001",
    "1111001100010001",
    "1111000110111110",
    "1111000000101100",
    "1110111001111010",
    "1110110011010101",
    "1110101101110000",
    "1110101001101101",
    "1110100111011011",
    "1110100110101010",
    "1110100110111110",
    "1110100111110001",
    "1110101000101000",
    "1110101001011011",
    "1110101001111101",
    "1110101010010100",
    "1110101010011110",
    "1110101010100101",
    "1110101010110101",
    "1110101011100101",
    "1110101101010001",
    "1110110000100001",
    "1110110101111001",
    "1110111101110010",
    "1111001000000100",
    "1111010100001010",
    "1111100001000000",
    "1111101101011000",
    "1111111000000110",
    "1111111111011100",
    "1111111001010011",
    "1111110100110010",
    "1111110000111011",
    "1111101100110100",
    "1111100111110110",
    "1111100010000000",
    "1111011011100101",
    "1111010101001110",
    "1111001111011110",
    "1111001010110000",
    "1111000111001001",
    "1111000100101001",
    "1111000011000011",
    "1111000010010111",
    "1111000010011101",
    "1111000011010000",
    "1111000100011100",
    "1111000101100000",
    "1111000101111100",
    "1111000101001101",
    "1111000010111110",
    "1110111111010111",
    "1110111010101101",
    "1110110101100111",
    "1110110000110011",
    "1110101100110000",
    "1110101001110101",
    "1110101000001011",
    "1110100111101100",
    "1110101000010000",
    "1110101001100011",
    "1110101011010100",
    "1110101101001110",
    "1110101110111111",
    "1110110000011100",
    "1110110001100110",
    "1110110010101001",
    "1110110011111001",
    "1110110101101100",
    "1110111000010110",
    "1110111100000001",
    "1111000000110000",
    "1111000110100010",
    "1111001101001110",
    "1111010100101100",
    "1111011100110101",
    "1111100101011010",
    "1111101110001100",
    "1111110110110010",
    "1111111110110100",
    "1111111010000110",
    "1111110100011001",
    "1111110000010001",
    "1111101101110101",
    "1111101101000101",
    "1111101101111001",
    "1111101111111111",
    "1111110010111010",
    "1111110110001011",
    "1111111001010000",
    "1111111011101010",
    "1111111101000001",
    "1111111101001000",
    "1111111011111010",
    "1111111001011111",
    "1111110110000101",
    "1111110001111110",
    "1111101101100000",
    "1111101000111001",
    "1111100100011101",
    "1111100000011001",
    "1111011101000000",
    "1111011010101010",
    "1111011001011101",
    "1111011001010101",
    "1111011001110010",
    "1111011001111111",
    "1111011001001001",
    "1111010110101000",
    "1111010010010101",
    "1111001100100110",
    "1111000110001101",
    "1110111111110011",
    "1110111001111010",
    "1110110100110110",
    "1110110000100100",
    "1110101101000010",
    "1110101010001001",
    "1110100111110111",
    "1110100110001110",
    "1110100101001001",
    "1110100100100100",
    "1110100100010011",
    "1110100100001011",
    "1110100100001000",
    "1110100100000001",
    "1110100100000000",
    "1110100100010010",
    "1110100101001110",
    "1110100111001110",
    "1110101010100011",
    "1110101111000101",
    "1110110100011101",
    "1110111010000100",
    "1110111111011110",
    "1111000100011100",
    "1111001001000001",
    "1111001101010111",
    "1111010001100010",
    "1111010101010111",
    "1111011000011000",
    "1111011010000111",
    "1111011010010100",
    "1111011001000110",
    "1111010110110100",
    "1111010100000011",
    "1111010001010010",
    "1111001110110011",
    "1111001100101010",
    "1111001010110000",
    "1111001001000110",
    "1111000111110001",
    "1111000110111110",
    "1111000111000011",
    "1111001000001000",
    "1111001010001100",
    "1111001101000000",
    "1111010000000111",
    "1111010010111110",
    "1111010101001011",
    "1111010110011000",
    "1111010110011101",
    "1111010101011000",
    "1111010011011010",
    "1111010000110110",
    "1111001110001010",
    "1111001011110011",
    "1111001010001001",
    "1111001001011101",
    "1111001001110111",
    "1111001011001111",
    "1111001101011100",
    "1111010000001010",
    "1111010011001011",
    "1111010110011011",
    "1111011001111010",
    "1111011101101001",
    "1111100001100111",
    "1111100101101111",
    "1111101001101111",
    "1111101101010000",
    "1111101111110111",
    "1111110001010000",
    "1111110001010010",
    "1111101111111100",
    "1111101101011001",
    "1111101001111000",
    "1111100101101010",
    "1111100001000011",
    "1111011100010111",
    "1111011000000011",
    "1111010100100111",
    "1111010010100001",
    "1111010001111110",
    "1111010010111001",
    "1111010100110100",
    "1111010111001001",
    "1111011001011101",
    "1111011011100101",
    "1111011101101011",
    "1111100000000101",
    "1111100011001011",
    "1111100111000101",
    "1111101011101100",
    "1111110000101110",
    "1111110101110111",
    "1111111010111111",
    "1111111111111000",
    "1111111010101100",
    "1111110101010111",
    "1111101111111001",
    "1111101010011100",
    "1111100101010000",
    "1111100000100100",
    "1111011100101101",
    "1111011001111010",
    "1111011000011101",
    "1111011000100111",
    "1111011010100011",
    "1111011110010010",
    "1111100011101100",
    "1111101010011001",
    "1111110001111010",
    "1111111001101111",
    "1111111110100100",
    "1111110111100010",
    "1111110001100010",
    "1111101100110100",
    "1111101001011110",
    "1111100111011011",
    "1111100110101011",
    "1111100111001100",
    "1111101001000000",
    "1111101100001110",
    "1111110000110111",
    "1111110110101110",
    "1111111101011010",
    "1111111011100100",
    "1111110100110110",
    "1111101110111000",
    "1111101010000000",
    "1111100110011100",
    "1111100100001101",
    "1111100011001010",
    "1111100010111011",
    "1111100011000101",
    "1111100011000011",
    "1111100010010101",
    "1111100000110101",
    "1111011110101001",
    "1111011100010011",
    "1111011010011011",
    "1111011001100000",
    "1111011001110111",
    "1111011011011011",
    "1111011101111101",
    "1111100001000011",
    "1111100100011101",
    "1111101000000011",
    "1111101011110100",
    "1111101111110101",
    "1111110011111110",
    "1111110111111100",
    "1111111011001101",
    "1111111101001100",
    "1111111101010100",
    "1111111011010000",
    "1111110111000010",
    "1111110001001011",
    "1111101010100101",
    "1111100100010111",
    "1111011111101001",
    "1111011101010111",
    "1111011110001001",
    "1111100010000101",
    "1111101000101100",
    "1111110000111100",
    "1111111001100000",
    "1111111111000010",
    "1111111001111110",
    "1111111000000000",
    "1111111001001101",
    "1111111101000101",
    "1111111101010000",
    "1111110110110011",
    "1111110000011011",
    "1111101010101000",
    "1111100101101100",
    "1111100001100111",
    "1111011110001101",
    "1111011011001111",
    "1111011000100010",
    "1111010110000100",
    "1111010100001011",
    "1111010011001111",
    "1111010011101010",
    "1111010101110001",
    "1111011001100111",
    "1111011110111111",
    "1111100101011111",
    "1111101100101101",
    "1111110100001011",
    "1111111011011110",
    "1111111101101111",
    "1111110111111110",
    "1111110011100110",
    "1111110000111110",
    "1111110000001111",
    "1111110001010101",
    "1111110011111110",
    "1111110111101111",
    "1111111100001000",
    "1111111111001010",
    "1111111010010111",
    "1111110101010000",
    "1111101111100010",
    "1111101000111001",
    "1111100001000111",
    "1111011000001000",
    "1111001110000010",
    "1111000010111110",
    "1110110111010000",
    "1110101011010100",
    "1110011111111000",
    "1110010101101110",
    "1110001101011100",
    "1110000111011111",
    "1110000011110110",
    "1110000010001000",
    "1110000001110000",
    "1110000010001010",
    "1110000011000101",
    "1110000100100000",
    "1110000110101010",
    "1110001001111100",
    "1110001110110011",
    "1110010101101100",
    "1110011110110011",
    "1110101010000110",
    "1110110111001101",
    "1111000101011101",
    "1111010100000101",
    "1111100010010000",
    "1111101111001110",
    "1111111010011001",
    "1111111100101100",
    "1111110110010011",
    "1111110010001110",
    "1111110000000101",
    "1111101111001110",
    "1111101110111100",
    "1111101110101010",
    "1111101110000011",
    "1111101101001010",
    "1111101100011000",
    "1111101100010001",
    "1111101101011001",
    "1111110000000111",
    "1111110100100001",
    "1111111010011100",
    "1111111110100001",
    "1111110110111101",
    "1111101111011100",
    "1111101000101001",
    "1111100011010010",
    "1111100000000010",
    "1111011111011110",
    "1111100001111000",
    "1111100111000101",
    "1111101110011110",
    "1111110111001100",
    "1111111111110100",
    "1111110111100010",
    "1111110000100111",
    "1111101011010011",
    "1111100111011111",
    "1111100100101111",
    "1111100010100100",
    "1111100000100011",
    "1111011110011011",
    "1111011100001111",
    "1111011010001001",
    "1111011000011000",
    "1111010111000100",
    "1111010110001110",
    "1111010101101111",
    "1111010101100010",
    "1111010101011011",
    "1111010101010111",
    "1111010101010010",
    "1111010101001110",
    "1111010101010011",
    "1111010101100000",
    "1111010101111110",
    "1111010110101100",
    "1111010111101000",
    "1111011000110010",
    "1111011010000100",
    "1111011011010110",
    "1111011100100110",
    "1111011101110000",
    "1111011110111010",
    "1111100000001101",
    "1111100001111000",
    "1111100100000101",
    "1111100110111100",
    "1111101010100111",
    "1111101111010001",
    "1111110101000111",
    "1111111100010110",
    "1111111010111000",
    "1111110000110001",
    "1111100101110010",
    "1111011010110010",
    "1111010000101001",
    "1111001000001011",
    "1111000001101110",
    "1110111101001001",
    "1110111001110101",
    "1110110111000011",
    "1110110100001011",
    "1110110001000010",
    "1110101101101011",
    "1110101010100010",
    "1110100111110111",
    "1110100101110001",
    "1110100100001000",
    "1110100010100111",
    "1110100000111101",
    "1110011111000111",
    "1110011101010010",
    "1110011011111000",
    "1110011011010110",
    "1110011011111100",
    "1110011101100110",
    "1110011111111011",
    "1110100010010010",
    "1110100100000011",
    "1110100100111001",
    "1110100100110001",
    "1110100100000101",
    "1110100011010111",
    "1110100011010011",
    "1110100100011010",
    "1110100110111100",
    "1110101010111111",
    "1110110000011001",
    "1110110110110111",
    "1110111110000101",
    "1111000101101100",
    "1111001101001111",
    "1111010100010010",
    "1111011010010001",
    "1111011110110000",
    "1111100001011100",
    "1111100010010111",
    "1111100001110110",
    "1111100000011100",
    "1111011110110110",
    "1111011101110010",
    "1111011101101110",
    "1111011110111011",
    "1111100001011010",
    "1111100100111100",
    "1111101001000110",
    "1111101101100000",
    "1111110001111001",
    "1111110110001001",
    "1111111010010010",
    "1111111110010111",
    "1111111101101000",
    "1111111001110110",
    "1111110110011100",
    "1111110011011001",
    "1111110000100100",
    "1111101101100110",
    "1111101010001000",
    "1111100101101111",
    "1111100000001100",
    "1111011001010001",
    "1111010000111011",
    "1111000111000100",
    "1110111011110101",
    "1110101111011110",
    "1110100010100001",
    "1110010101101010",
    "1110001001101011",
    "1101111111010001",
    "1101110110111111",
    "1101110001001101",
    "1101101110000101",
    "1101101101101001",
    "1101101111111010",
    "1101110100101001",
    "1101111011100101",
    "1110000100010000",
    "1110001110000100",
    "1110011000011110",
    "1110100011000011",
    "1110101101100000",
    "1110110111101000",
    "1111000001010000",
    "1111001010000111",
    "1111010001111001",
    "1111011000010101",
    "1111011101010001",
    "1111100000110110",
    "1111100011011010",
    "1111100101011000",
    "1111100111001010",
    "1111101000111100",
    "1111101010101111",
    "1111101100010111",
    "1111101101100111",
    "1111101110010011",
    "1111101110011011",
    "1111101110001010",
    "1111101101111000",
    "1111101101111111",
    "1111101110101101",
    "1111110000000011",
    "1111110001101111",
    "1111110011010010",
    "1111110100001011",
    "1111110011111101",
    "1111110010011111",
    "1111101111110010",
    "1111101100000111",
    "1111100111110100",
    "1111100011001000",
    "1111011110001111",
    "1111011001001100",
    "1111010011111000",
    "1111001110000000",
    "1111000111010110",
    "1110111111110011",
    "1110110111101010",
    "1110101111100110",
    "1110101000100000",
    "1110100011010000",
    "1110100000100001",
    "1110100000011110",
    "1110100010111001",
    "1110100111001110",
    "1110101100111000",
    "1110110011010011",
    "1110111010001100",
    "1111000001010101",
    "1111001000100000",
    "1111001111011001",
    "1111010101100100",
    "1111011010100101",
    "1111011110000100",
    "1111011111110001",
    "1111011111101110",
    "1111011110001010",
    "1111011011011011",
    "1111010111110101",
    "1111010011101001",
    "1111001111000100",
    "1111001010001111",
    "1111000101100000",
    "1111000001001000",
    "1110111101011011",
    "1110111010101000",
    "1110111000110111",
    "1110111000001110",
    "1110111000101010",
    "1110111010000110",
    "1110111100011110",
    "1110111111101001",
    "1111000011010111",
    "1111000111010101",
    "1111001011010100",
    "1111001111001000",
    "1111010010110100",
    "1111010110100000",
    "1111011010010100",
    "1111011110011110",
    "1111100010111110",
    "1111100111110100",
    "1111101100110100",
    "1111110001110000",
    "1111110110011111",
    "1111111011000000",
    "1111111111001110",
    "1111111100110010",
    "1111111001001011",
    "1111110101111110",
    "1111110011011010",
    "1111110001110000",
    "1111110001010111",
    "1111110010101101",
    "1111110110001110",
    "1111111100011000",
    "1111111010100111",
    "1111101111001001",
    "1111100010001011",
    "1111010101010010",
    "1111001010001111",
    "1111000010100001",
    "1110111110110110",
    "1110111111000010",
    "1111000010001000",
    "1111000110110100",
    "1111001011110111",
    "1111010000011111",
    "1111010100011111",
    "1111010111111010",
    "1111011011000111",
    "1111011110010110",
    "1111100001110000",
    "1111100101010101",
    "1111101001000111",
    "1111101101000011",
    "1111110001001000",
    "1111110101011001",
    "1111111001110000",
    "1111111101111101",
    "1111111110010110",
    "1111111011101101",
    "1111111010011001",
    "1111111010011111",
    "1111111011110011",
    "1111111101110111",
    "1111111111110011",
    "1111111101110000",
    "1111111100001101",
    "1111111011010001",
    "1111111010110010",
    "1111111010100100",
    "1111111010011101",
    "1111111010010010",
    "1111111010000000",
    "1111111001101011",
    "1111111001011000",
    "1111111001001110",
    "1111111001010011",
    "1111111001101001",
    "1111111010001111",
    "1111111010111110",
    "1111111011100111",
    "1111111011111110",
    "1111111011110100",
    "1111111011000110",
    "1111111001110110",
    "1111111000010011",
    "1111110110101000",
    "1111110101000101",
    "1111110011110110",
    "1111110011000110",
    "1111110011000001",
    "1111110011110001",
    "1111110101100000",
    "1111111000010010",
    "1111111100000100",
    "1111111111010000",
    "1111111010000011",
    "1111110100100011",
    "1111101110111111",
    "1111101001011101",
    "1111100100000000",
    "1111011110100110",
    "1111011001010011",
    "1111010100001011",
    "1111001111011010",
    "1111001011010100",
    "1111001000001001",
    "1111000110001000",
    "1111000101100000",
    "1111000110011010",
    "1111001000110101",
    "1111001100100110",
    "1111010001010111",
    "1111010110100100",
    "1111011011100101",
    "1111011111110110",
    "1111100010110100",
    "1111100100001101",
    "1111100011111011",
    "1111100010001111",
    "1111011111101001",
    "1111011100110101",
    "1111011010011001",
    "1111011000110100",
    "1111011000001100",
    "1111011000011000",
    "1111011000111010",
    "1111011001010011",
    "1111011001000010",
    "1111010111110001",
    "1111010101001110",
    "1111010001010100",
    "1111001011111010",
    "1111000101000101",
    "1110111100111000",
    "1110110011100110",
    "1110101001100011",
    "1110011111001101",
    "1110010101001001",
    "1110001011110011",
    "1110000011100110",
    "1101111100101101",
    "1101110111010000",
    "1101110011001000",
    "1101110000001100",
    "1101101110010001",
    "1101101101001010",
    "1101101100110000",
    "1101101101000000",
    "1101101101111000",
    "1101101111011001",
    "1101110001100110",
    "1101110100100100",
    "1101111000100000",
    "1101111101101001",
    "1110000100011000",
    "1110001100111100",
    "1110010111011000",
    "1110100011011000",
    "1110110000010100",
    "1110111101010001",
    "1111001001010101",
    "1111010011101110",
    "1111011011110101",
    "1111100001011110",
    "1111100100101111",
    "1111100110000000",
    "1111100101111110",
    "1111100101100010",
    "1111100101101100",
    "1111100111011000",
    "1111101011001111",
    "1111110001011100",
    "1111111001101000",
    "1111111100111011",
    "1111110011010011",
    "1111101010011000",
    "1111100010110011",
    "1111011100101110",
    "1111011000000110",
    "1111010100100100",
    "1111010001110110",
    "1111001111110110",
    "1111001110101001",
    "1111001110010110",
    "1111001111000000",
    "1111010000100011",
    "1111010010111001",
    "1111010101111011",
    "1111011001100000",
    "1111011101101001",
    "1111100010010100",
    "1111100111011000",
    "1111101100100110",
    "1111110001011111",
    "1111110101011111",
    "1111111000000111",
    "1111111001001000",
    "1111111000101010",
    "1111110111001101",
    "1111110101011011",
    "1111110011111101",
    "1111110011010000",
    "1111110011011100",
    "1111110100010111",
    "1111110101101101",
    "1111110111000101",
    "1111111000001101",
    "1111111000110111",
    "1111111001000010",
    "1111111000110101",
    "1111111000011100",
    "1111111000000100",
    "1111110111110110",
    "1111110111111100",
    "1111111000011001",
    "1111111001001100",
    "1111111010001100",
    "1111111011000010",
    "1111111011010111",
    "1111111010110111",
    "1111111001011010",
    "1111110111001101",
    "1111110100101100",
    "1111110010101001",
    "1111110001110100",
    "1111110011000100",
    "1111110111001010",
    "1111111110101100",
    "1111110110000100",
    "1111100111101011",
    "1111010111010001",
    "1111000110101000",
    "1110110111100111",
    "1110101011110000",
    "1110100011111001",
    "1110100000000010",
    "1110011111100001",
    "1110100001011001",
    "1110100100100000",
    "1110100111111110",
    "1110101011000111",
    "1110101101100001",
    "1110101110111111",
    "1110101111011110",
    "1110101111000111",
    "1110101110001100",
    "1110101101000100",
    "1110101100000100",
    "1110101011100011",
    "1110101011101000",
    "1110101100010111",
    "1110101101101110",
    "1110101111100100",
    "1110110001110100",
    "1110110100011101",
    "1110110111011111",
    "1110111010111010",
    "1110111110101011",
    "1111000010101011",
    "1111000110110001",
    "1111001010101101",
    "1111001110010100",
    "1111010001010101",
    "1111010011100110",
    "1111010100111001",
    "1111010101010000",
    "1111010100101110",
    "1111010011011111",
    "1111010001111000",
    "1111010000001101",
    "1111001110111010",
    "1111001110001101",
    "1111001110010110",
    "1111001111010100",
    "1111010001000101",
    "1111010011100110",
    "1111010110101111",
    "1111011010100011",
    "1111011111000010",
    "1111100100001101",
    "1111101010000101",
    "1111110000101100",
    "1111111000000101",
    "1111111111101101",
    "1111110110101111",
    "1111101100111111",
    "1111100010100001",
    "1111010111100011",
    "1111001100011011",
    "1111000001110000",
    "1110111000010001",
    "1110110000110000",
    "1110101011101111",
    "1110101001011110",
    "1110101001110100",
    "1110101100001111",
    "1110110000000011",
    "1110110100100101",
    "1110111001010011",
    "1110111101101101",
    "1111000001100001",
    "1111000100011000",
    "1111000110000001",
    "1111000110001110",
    "1111000100111011",
    "1111000010010000",
    "1110111110100100",
    "1110111010010011",
    "1110110101111001",
    "1110110001100110",
    "1110101101100100",
    "1110101001101111",
    "1110100110000000",
    "1110100010010101",
    "1110011110111010",
    "1110011011111000",
    "1110011001101000",
    "1110011000011000",
    "1110011000010110",
    "1110011001100111",
    "1110011100001001",
    "1110011111110110",
    "1110100100011101",
    "1110101001101010",
    "1110101111000000",
    "1110110100000110",
    "1110111000100010",
    "1110111100000111",
    "1110111110101110",
    "1111000000011001",
    "1111000001001100",
    "1111000001010101",
    "1111000001000111",
    "1111000000111001",
    "1111000001001000",
    "1111000010000110",
    "1111000100000000",
    "1111000110101100",
    "1111001001110100",
    "1111001100110111",
    "1111001111011001",
    "1111010001000111",
    "1111010010000000",
    "1111010010001011",
    "1111010001110001",
    "1111010000111000",
    "1111001111011001",
    "1111001101001100",
    "1111001010000110",
    "1111000101111100",
    "1111000000110101",
    "1110111010110111",
    "1110110100100000",
    "1110101110010110",
    "1110101001000001",
    "1110100101001000",
    "1110100011001000",
    "1110100011010000",
    "1110100101011111",
    "1110101001100011",
    "1110101111000101",
    "1110110101101001",
    "1110111100110101",
    "1111000100010101",
    "1111001011110011",
    "1111010010111101",
    "1111011001100000",
    "1111011111001111",
    "1111100100000110",
    "1111101000000010",
    "1111101011001001",
    "1111101101100010",
    "1111101111001110",
    "1111110000001010",
    "1111110000010010",
    "1111101111011101",
    "1111101101101111",
    "1111101011010011",
    "1111101000011000",
    "1111100101010000",
    "1111100010000110",
    "1111011110111111",
    "1111011011101101",
    "1111011000001011",
    "1111010100001011",
    "1111001111110000",
    "1111001011000100",
    "1111000110100100",
    "1111000010110011",
    "1111000000011100",
    "1110111111111111",
    "1111000001110011",
    "1111000101111001",
    "1111001011111101",
    "1111010011011101",
    "1111011011110101",
    "1111100100011000",
    "1111101100100100",
    "1111110100000001",
    "1111111010011101",
    "1111111111110001",
    "1111111100000000",
    "1111111000110100",
    "1111110110100000",
    "1111110100111110",
    "1111110100001001",
    "1111110011111100",
    "1111110100010000",
    "1111110100110111",
    "1111110101011110",
    "1111110101110101",
    "1111110101110101",
    "1111110101100110",
    "1111110101100001",
    "1111110110000010",
    "1111110111100101",
    "1111111010011011",
    "1111111110101100",
    "1111111011101100",
    "1111110101000001",
    "1111101101100111",
    "1111100101111011",
    "1111011110011100",
    "1111010111101101",
    "1111010010001011",
    "1111001110000010",
    "1111001011010100",
    "1111001001110100",
    "1111001001010001",
    "1111001001100000",
    "1111001010011101",
    "1111001100000111",
    "1111001110101101",
    "1111010010010111",
    "1111010111001101",
    "1111011101001111",
    "1111100100011100",
    "1111101100101110",
    "1111110101111001",
    "1111111111101011",
    "1111110110010001",
    "1111101100100000",
    "1111100011011100",
    "1111011011100001",
    "1111010101000001",
    "1111010000000011",
    "1111001100011110",
    "1111001001111010",
    "1111000111111110",
    "1111000110001011",
    "1111000100010000",
    "1111000010000110",
    "1110111111111000",
    "1110111101111111",
    "1110111100111000",
    "1110111100111010",
    "1110111110010010",
    "1111000000111110",
    "1111000100101111",
    "1111001001010101",
    "1111001110010100",
    "1111010011011101",
    "1111011000011110",
    "1111011101001100",
    "1111100001011111",
    "1111100101010010",
    "1111101000100011",
    "1111101011010111",
    "1111101101110111",
    "1111110000000010",
    "1111110001110100",
    "1111110010111001",
    "1111110010111010",
    "1111110001100010",
    "1111101110100110",
    "1111101010001100",
    "1111100100101010",
    "1111011110100011",
    "1111011000010101",
    "1111010010010111",
    "1111001100110000",
    "1111000111010110",
    "1111000010000101",
    "1110111100111101",
    "1110111000010001",
    "1110110100100101",
    "1110110010100001",
    "1110110010101100",
    "1110110101011011",
    "1110111010110000",
    "1111000010011001",
    "1111001011111000",
    "1111010110100101",
    "1111100001101110",
    "1111101100011010",
    "1111110101110001",
    "1111111101001001",
    "1111111101110100",
    "1111111011001110",
    "1111111010110000",
    "1111111011111101",
    "1111111110010101",
    "1111111110011110",
    "1111111010110011",
    "1111110110101010",
    "1111110010000101",
    "1111101100111111",
    "1111100111011011",
    "1111100001010111",
    "1111011010110010",
    "1111010011100111",
    "1111001011110010",
    "1111000011001010",
    "1110111001101111",
    "1110101111101110",
    "1110100101011010",
    "1110011011010100",
    "1110010001111001",
    "1110001001100000",
    "1110000010010000",
    "1101111100010001",
    "1101110111011111",
    "1101110011111110",
    "1101110001111000",
    "1101110001011001",
    "1101110010110100",
    "1101110110010010",
    "1101111011110011",
    "1110000011010111",
    "1110001100111111",
    "1110011000110010",
    "1110100110110010",
    "1110110110111001",
    "1111001000100011",
    "1111011010110100",
    "1111101100011100",
    "1111111100010001",
    "1111110110100001",
    "1111101100011111",
    "1111100101100101",
    "1111100001011111",
    "1111011111101011",
    "1111011111100100",
    "1111100000101110",
    "1111100010101110",
    "1111100101011000",
    "1111101000100011",
    "1111101100010100",
    "1111110000110101",
    "1111110110010010",
    "1111111100110010",
    "1111111011110100",
    "1111110100001000",
    "1111101101000011",
    "1111100111101110",
    "1111100101010010",
    "1111100110011101",
    "1111101011010111",
    "1111110011011100",
    "1111111101100011",
    "1111110111101001",
    "1111101101100011",
    "1111100101000110",
    "1111011110110110",
    "1111011010110010",
    "1111011000011101",
    "1111010111001001",
    "1111010110000011",
    "1111010100100010",
    "1111010010001111",
    "1111001111000111",
    "1111001011011000",
    "1111000111011111",
    "1111000011111011",
    "1111000001001101",
    "1110111111101001",
    "1110111111011001",
    "1111000000010100",
    "1111000010010000",
    "1111000100110011",
    "1111000111100111",
    "1111001010011000",
    "1111001100111000",
    "1111001111000000",
    "1111010000101110",
    "1111010010000110",
    "1111010011010011",
    "1111010100011100",
    "1111010101100111",
    "1111010110111100",
    "1111011000011000",
    "1111011001110101",
    "1111011011001010",
    "1111011100001001",
    "1111011100101000",
    "1111011100100011",
    "1111011100000111",
    "1111011011110011",
    "1111011100010011",
    "1111011110010100",
    "1111100010011010",
    "1111101000101111",
    "1111110001000001",
    "1111111010100111",
    "1111111011001011",
    "1111110001010010",
    "1111101000010101",
    "1111100000110001",
    "1111011010110000",
    "1111010110001011",
    "1111010010101001",
    "1111001111100110",
    "1111001100010110",
    "1111001000010001",
    "1111000011000011",
    "1110111100101010",
    "1110110101011010",
    "1110101101111010",
    "1110100110110111",
    "1110100000110110",
    "1110011100000101",
    "1110011000100010",
    "1110010101111100",
    "1110010011111011",
    "1110010010001010",
    "1110010000100011",
    "1110001111000111",
    "1110001110000100",
    "1110001101100100",
    "1110001101111000",
    "1110001111001101",
    "1110010001110110",
    "1110010101111100",
    "1110011011101000",
    "1110100010110100",
    "1110101011010001",
    "1110110100011101",
    "1110111101110011",
    "1111000110101111",
    "1111001110101101",
    "1111010101010010",
    "1111011010001111",
    "1111011101100000",
    "1111011111000000",
    "1111011110111111",
    "1111011101101101",
    "1111011011100011",
    "1111011001000010",
    "1111010110101000",
    "1111010100101110",
    "1111010011100100",
    "1111010011001111",
    "1111010011101111",
    "1111010101000011",
    "1111010111000110",
    "1111011001110100",
    "1111011101000111",
    "1111100000111000",
    "1111100100110011",
    "1111101000100101",
    "1111101011111001",
    "1111101110100000",
    "1111110000011101",
    "1111110010000000",
    "1111110011101001",
    "1111110101111101",
    "1111111001010111",
    "1111111110001011",
    "1111111011101000",
    "1111110100010110",
    "1111101100001001",
    "1111100011001011",
    "1111011001011110",
    "1111001110111111",
    "1111000011101001",
    "1110110111100111",
    "1110101011001001",
    "1110011110110001",
    "1110010010111110",
    "1110001000001100",
    "1101111110110011",
    "1101110110111111",
    "1101110000111001",
    "1101101100100110",
    "1101101010001111",
    "1101101001111100",
    "1101101011111100",
    "1101110000010101",
    "1101110111001011",
    "1110000000001101",
    "1110001010110111",
    "1110010110010110",
    "1110100001111000",
    "1110101100110101",
    "1110110110111001",
    "1111000000000101",
    "1111001000100010",
    "1111010000011001",
    "1111010111101000",
    "1111011110000101",
    "1111100011100001",
    "1111100111110001",
    "1111101010111001",
    "1111101101001000",
    "1111101110110010",
    "1111110000001110",
    "1111110001110000",
    "1111110011100110",
    "1111110101111001",
    "1111111000101001",
    "1111111011101101",
    "1111111110110110",
    "1111111110001011",
    "1111111011110001",
    "1111111010001010",
    "1111111001100010",
    "1111111001111101",
    "1111111011011011",
    "1111111101111011",
    "1111111110100000",
    "1111111001111010",
    "1111110100001100",
    "1111101101010110",
    "1111100101011011",
    "1111011100100110",
    "1111010011001010",
    "1111001001100011",
    "1111000000011100",
    "1110111000110000",
    "1110110011010101",
    "1110110000110011",
    "1110110001011010",
    "1110110100110110",
    "1110111010011000",
    "1111000001000000",
    "1111000111101101",
    "1111001101110010",
    "1111010010101111",
    "1111010110100100",
    "1111011001011000",
    "1111011011100000",
    "1111011101001111",
    "1111011110110110",
    "1111100000011001",
    "1111100001110000",
    "1111100010101110",
    "1111100010111110",
    "1111100010001010",
    "1111100000000010",
    "1111011100100001",
    "1111010111101101",
    "1111010001111000",
    "1111001011011101",
    "1111000100110100",
    "1110111110011111",
    "1110111000111001",
    "1110110100011010",
    "1110110001010111",
    "1110101111111101",
    "1110110000001100",
    "1110110001111000",
    "1110110100101110",
    "1110111000010110",
    "1110111100100000",
    "1111000000111101",
    "1111000101101010",
    "1111001010110010",
    "1111010000011111",
    "1111010110111100",
    "1111011110001001",
    "1111100101111011",
    "1111101110000011",
    "1111110110000101",
    "1111111101100000",
    "1111111100001010",
    "1111110111010111",
    "1111110100010011",
    "1111110010111101",
    "1111110011000011",
    "1111110100001011",
    "1111110101111000",
    "1111110111110111",
    "1111111010000110",
    "1111111100110011",
    "1111111111100100",
    "1111111010101011",
    "1111110100010000",
    "1111101100100000",
    "1111100100000000",
    "1111011011100110",
    "1111010100010101",
    "1111001110111010",
    "1111001011101111",
    "1111001010101101",
    "1111001011100000",
    "1111001101100100",
    "1111010000011111",
    "1111010011111011",
    "1111010111110100",
    "1111011100000100",
    "1111100000101011",
    "1111100101100101",
    "1111101010101010",
    "1111101111101110",
    "1111110100101110",
    "1111111001110001",
    "1111111110111101",
    "1111111011100011",
    "1111110101111011",
    "1111110000100011",
    "1111101100000110",
    "1111101001010101",
    "1111101000111000",
    "1111101010111011",
    "1111101111001101",
    "1111110100111101",
    "1111111011001001",
    "1111111111001100",
    "1111111010111011",
    "1111111000010011",
    "1111110111001101",
    "1111110111001100",
    "1111110111101101",
    "1111111000010011",
    "1111111000101011",
    "1111111000101100",
    "1111111000011010",
    "1111110111111011",
    "1111110111010110",
    "1111110110110000",
    "1111110110001100",
    "1111110101101110",
    "1111110101010100",
    "1111110101000000",
    "1111110100110101",
    "1111110100110111",
    "1111110101001110",
    "1111110101111110",
    "1111110111001010",
    "1111111000110010",
    "1111111010110101",
    "1111111101001100",
    "1111111111110110",
    "1111111101010001",
    "1111111010010010",
    "1111110111010010",
    "1111110100010110",
    "1111110001011100",
    "1111101110100001",
    "1111101011011011",
    "1111100111111001",
    "1111100011110100",
    "1111011111000111",
    "1111011001110000",
    "1111010100000000",
    "1111001110000111",
    "1111001000100011",
    "1111000011110100",
    "1111000000011110",
    "1110111110110000",
    "1110111110110000",
    "1111000000010001",
    "1111000010111001",
    "1111000110001110",
    "1111001001111010",
    "1111001101110000",
    "1111010001101011",
    "1111010101100010",
    "1111011001000110",
    "1111011100000001",
    "1111011101111101",
    "1111011110101001",
    "1111011110000101",
    "1111011100100000",
    "1111011010011001",
    "1111011000010011",
    "1111010110101000",
    "1111010101101111",
    "1111010101101001",
    "1111010110001101",
    "1111010111001011",
    "1111011000010000",
    "1111011000111111",
    "1111011001000010",
    "1111010111111010",
    "1111010101001110",
    "1111010000100111",
    "1111001001111111",
    "1111000001100110",
    "1110111000001001",
    "1110101110100110",
    "1110100110000000",
    "1110011111001100",
    "1110011010100010",
    "1110010111110101",
    "1110010110011010",
    "1110010101010111",
    "1110010011111110",
    "1110010001111011",
    "1110001111010100",
    "1110001100101011",
    "1110001010101011",
    "1110001001111100",
    "1110001010111000",
    "1110001101100100",
    "1110010001110000",
    "1110010110111001",
    "1110011100010111",
    "1110100001101100",
    "1110100110100101",
    "1110101011000001",
    "1110101111010100",
    "1110110100000011",
    "1110111001101101",
    "1111000000100001",
    "1111001000011010",
    "1111010000110101",
    "1111011001000001",
    "1111100000001010",
    "1111100101101110",
    "1111101001100001",
    "1111101011111100",
    "1111101101110000",
    "1111101111111000",
    "1111110011001110",
    "1111111000010100",
    "1111111111010010",
    "1111111000001100",
    "1111101110111011",
    "1111100101101110",
    "1111011101010010",
    "1111010110001011",
    "1111010000100100",
    "1111001100011110",
    "1111001001101101",
    "1111001000000100",
    "1111000111011000",
    "1111000111100000",
    "1111001000010101",
    "1111001001110000",
    "1111001011110000",
    "1111001110001111",
    "1111010001001000",
    "1111010100011100",
    "1111010111111010",
    "1111011011100000",
    "1111011110111000",
    "1111100001111001",
    "1111100100011010",
    "1111100110010101",
    "1111100111101100",
    "1111101000100111",
    "1111101001010101",
    "1111101010000000",
    "1111101010110010",
    "1111101011101100",
    "1111101100101001",
    "1111101101100010",
    "1111101110001110",
    "1111101110101010",
    "1111101110110111",
    "1111101110111011",
    "1111101110111101",
    "1111101111000110",
    "1111101111011000",
    "1111101111110101",
    "1111110000011011",
    "1111110001001000",
    "1111110001110010",
    "1111110010001111",
    "1111110010001111",
    "1111110001101001",
    "1111110000010110",
    "1111101110100001",
    "1111101100011110",
    "1111101010101011",
    "1111101001101001",
    "1111101001110010",
    "1111101011011001",
    "1111101110100110",
    "1111110011011010",
    "1111111001110001",
    "1111111110010110",
    "1111110101000110",
    "1111101010100000",
    "1111011110110101",
    "1111010010100110",
    "1111000110100000",
    "1110111011100001",
    "1110110010011100",
    "1110101011110000",
    "1110100111100101",
    "1110100101100101",
    "1110100101000011",
    "1110100101010101",
    "1110100101110111",
    "1110100110010011",
    "1110100110100111",
    "1110100110110010",
    "1110100110111011",
    "1110100111000110",
    "1110100111010011",
    "1110100111100111",
    "1110101000000110",
    "1110101000110111",
    "1110101010000110",
    "1110101011111100",
    "1110101110011011",
    "1110110001011111",
    "1110110101000000",
    "1110111000110100",
    "1110111100111000",
    "1111000001001010",
    "1111000101100101",
    "1111001001111101",
    "1111001110000010",
    "1111010001011110",
    "1111010011110100",
    "1111010100110110",
    "1111010100010111",
    "1111010010011001",
    "1111001111010010",
    "1111001011100000",
    "1111000111101100",
    "1111000100100010",
    "1111000010100111",
    "1111000010010101",
    "1111000011110100",
    "1111000110111100",
    "1111001011011001",
    "1111010000110011",
    "1111010110110001",
    "1111011101000100",
    "1111100011100110",
    "1111101010100001",
    "1111110001111111",
    "1111111010001010",
    "1111111100111000",
    "1111110011010111",
    "1111101001100100",
    "1111100000000010",
    "1111010111011011",
    "1111010000011100",
    "1111001011100001",
    "1111001000111010",
    "1111001000011101",
    "1111001001101011",
    "1111001011111010",
    "1111001110011100",
    "1111010000110001",
    "1111010010100110",
    "1111010011111000",
    "1111010100101111",
    "1111010101010101",
    "1111010101101110",
    "1111010101110001",
    "1111010101001110",
    "1111010011111011",
    "1111010001100111",
    "1111001110010110",
    "1111001010010001",
    "1111000101101001",
    "1111000000110110",
    "1110111100010001",
    "1110111000010001",
    "1110110101000110",
    "1110110010110001",
    "1110110001000000",
    "1110101111010010",
    "1110101101000000",
    "1110101001101101",
    "1110100101010011",
    "1110100000000111",
    "1110011010110111",
    "1110010110011101",
    "1110010011101100",
    "1110010011000001",
    "1110010100100010",
    "1110010111111001",
    "1110011100100011",
    "1110100001111110",
    "1110100111110100",
    "1110101101111010",
    "1110110100010011",
    "1110111011000111",
    "1111000010011010",
    "1111001001111001",
    "1111010001001010",
    "1111010111101000",
    "1111011100110000",
    "1111100000001010",
    "1111100001110001",
    "1111100001110001",
    "1111100000100110",
    "1111011110110101",
    "1111011101000010",
    "1111011011101011",
    "1111011010111101",
    "1111011010111100",
    "1111011011010001",
    "1111011011011101",
    "1111011010110101",
    "1111011000110000",
    "1111010100110110",
    "1111001110111101",
    "1111000111100010",
    "1110111111011100",
    "1110110111110001",
    "1110110001101011",
    "1110101101111000",
    "1110101100101110",
    "1110101101111101",
    "1110110000111110",
    "1110110101001001",
    "1110111010000010",
    "1110111111011110",
    "1111000101011011",
    "1111001011111101",
    "1111010010111001",
    "1111011001110111",
    "1111100000011001",
    "1111100101110111",
    "1111101001111011",
    "1111101100010101",
    "1111101101001000",
    "1111101100100001",
    "1111101010110111",
    "1111101000100101",
    "1111100110000100",
    "1111100011101110",
    "1111100001110001",
    "1111100000010100",
    "1111011111001111",
    "1111011110010110",
    "1111011101000111",
    "1111011011000010",
    "1111010111100101",
    "1111010010100001",
    "1111001100000100",
    "1111000100111001",
    "1110111110000100",
    "1110111000101111",
    "1110110101111011",
    "1110110110000110",
    "1110111001001011",
    "1110111110100011",
    "1111000101010111",
    "1111001100101101",
    "1111010011110100",
    "1111011010001100",
    "1111011111101011",
    "1111100100010101",
    "1111101000011000",
    "1111101100000011",
    "1111101111100100",
    "1111110011000010",
    "1111110110010110",
    "1111111001010011",
    "1111111011100101",
    "1111111100111101",
    "1111111101011011",
    "1111111101001101",
    "1111111100101110",
    "1111111100100011",
    "1111111101001000",
    "1111111110101101",
    "1111111110110010",
    "1111111011110110",
    "1111111001000010",
    "1111110111000100",
    "1111110110100111",
    "1111111000001010",
    "1111111011111101",
    "1111111110000100",
    "1111110110011001",
    "1111101101101000",
    "1111100100100010",
    "1111011011110000",
    "1111010011110100",
    "1111001101000100",
    "1111000111100111",
    "1111000011011000",
    "1111000000011001",
    "1110111110100110",
    "1110111110000111",
    "1110111111001000",
    "1111000001110011",
    "1111000110001110",
    "1111001100010110",
    "1111010011111100",
    "1111011100101101",
    "1111100110001001",
    "1111101111111001",
    "1111111001100100",
    "1111111101001000",
    "1111110100011110",
    "1111101100100011",
    "1111100101100000",
    "1111011111011110",
    "1111011010101010",
    "1111010111010101",
    "1111010101101110",
    "1111010101110110",
    "1111010111100010",
    "1111011010010110",
    "1111011101101101",
    "1111100000111001",
    "1111100011011000",
    "1111100100110110",
    "1111100101010000",
    "1111100100110001",
    "1111100011110100",
    "1111100010110110",
    "1111100010010000",
    "1111100010010100",
    "1111100011000101",
    "1111100100011100",
    "1111100110000110",
    "1111100111101011",
    "1111101000110001",
    "1111101001000001",
    "1111101000001111",
    "1111100110011000",
    "1111100011101001",
    "1111100000001101",
    "1111011100010111",
    "1111011000010110",
    "1111010100010010",
    "1111010000010111",
    "1111001100110000",
    "1111001001100101",
    "1111000110111100",
    "1111000100110110",
    "1111000011010000",
    "1111000010001101",
    "1111000001101100",
    "1111000001110000",
    "1111000010010101",
    "1111000011011000",
    "1111000100101111",
    "1111000110010011",
    "1111001000000011",
    "1111001010000111",
    "1111001100110101",
    "1111010000011111",
    "1111010101010010",
    "1111011011010001",
    "1111100010001101",
    "1111101001101001",
    "1111110000111110",
    "1111110111100011",
    "1111111100111011",
    "1111111111001100",
    "1111111100111011",
    "1111111100000011",
    "1111111100010111",
    "1111111101101010",
    "1111111111110011",
    "1111111101001001",
    "1111111001010101",
    "1111110100101101",
    "1111101111011010",
    "1111101001100000",
    "1111100010111110",
    "1111011011100110",
    "1111010011000110",
    "1111001001000110",
    "1110111101010010",
    "1110101111110110",
    "1110100001010101",
    "1110010010101111",
    "1110000101001011",
    "1101111001100011",
    "1101110000011010",
    "1101101001111101",
    "1101100101111100",
    "1101100100000101",
    "1101100100000001",
    "1101100101101111",
    "1101101001001001",
    "1101101110010001",
    "1101110100111110",
    "1101111101010001",
    "1110000111001101",
    "1110010010110100",
    "1110100000000101",
    "1110101110110000",
    "1110111110011100",
    "1111001110011111",
    "1111011110000100",
    "1111101100010110",
    "1111111000101000",
    "1111111101100001",
    "1111110110011100",
    "1111110010000101",
    "1111110000001110",
    "1111110000011101",
    "1111110010001111",
    "1111110101000001",
    "1111111000010011",
    "1111111011101110",
    "1111111111000110",
    "1111111101011110",
    "1111111001111100",
    "1111110110000100",
    "1111110001101111",
    "1111101101000111",
    "1111101000100100",
    "1111100100101111",
    "1111100010010111",
    "1111100010000110",
    "1111100100011100",
    "1111101001011000",
    "1111110000100101",
    "1111111001010011",
    "1111111101010111",
    "1111110100011100",
    "1111101100101001",
    "1111100110011111",
    "1111100010001010",
    "1111011111011100",
    "1111011110000000",
    "1111011101010110",
    "1111011100111100",
    "1111011100001111",
    "1111011010111101",
    "1111011000111010",
    "1111010110001011",
    "1111010011000001",
    "1111001111111011",
    "1111001101010100",
    "1111001011100101",
    "1111001010111100",
    "1111001011011001",
    "1111001100110000",
    "1111001110100110",
    "1111010000100100",
    "1111010010010111",
    "1111010011110001",
    "1111010100110100",
    "1111010101100111",
    "1111010110011000",
    "1111010111010101",
    "1111011000100000",
    "1111011001111111",
    "1111011011101000",
    "1111011101010001",
    "1111011110110000",
    "1111011111111000",
    "1111100000101001",
    "1111100001000101",
    "1111100001011111",
    "1111100010001010",
    "1111100011100010",
    "1111100101111001",
    "1111101001011000",
    "1111101101111110",
    "1111110011011011",
    "1111111001011101",
    "1111111111101110",
    "1111111001111101",
    "1111110011111110",
    "1111101110011101",
    "1111101001011111",
    "1111100101000101",
    "1111100001000010",
    "1111011101000000",
    "1111011000101010",
    "1111010011100100",
    "1111001101011100",
    "1111000110001101",
    "1110111110000010",
    "1110110101010011",
    "1110101100011100",
    "1110100100000001",
    "1110011100100011",
    "1110010110011011",
    "1110010001111000",
    "1110001110111101",
    "1110001101100011",
    "1110001101011100",
    "1110001110011001",
    "1110010000001101",
    "1110010010110011",
    "1110010110011010",
    "1110011011010001",
    "1110100001100100",
    "1110101001000111",
    "1110110001011100",
    "1110111001101101",
    "1111000001000011",
    "1111000110110100",
    "1111001010110000",
    "1111001101000000",
    "1111001110001001",
    "1111001110101110",
    "1111001111010100",
    "1111010000001010",
    "1111010001010111",
    "1111010010111000",
    "1111010100100100",
    "1111010110011010",
    "1111011000011101",
    "1111011010101111",
    "1111011101001010",
    "1111011111101000",
    "1111100001110100",
    "1111100011100010",
    "1111100100101100",
    "1111100101011011",
    "1111100101111100",
    "1111100110011011",
    "1111100110111110",
    "1111100111100011",
    "1111101000000110",
    "1111101000100011",
    "1111101001000001",
    "1111101001101010",
    "1111101010110000",
    "1111101100100011",
    "1111101111010100",
    "1111110011001011",
    "1111111000010110",
    "1111111111000010",
    "1111111000100001",
    "1111101110001010",
    "1111100001101001",
    "1111010011000000",
    "1111000010101011",
    "1110110001011111",
    "1110100000110001",
    "1110010001111000",
    "1110000101111110",
    "1101111101101000",
    "1101111000101111",
    "1101110110101010",
    "1101110110011000",
    "1101110110111100",
    "1101110111110010",
    "1101111000110101",
    "1101111010011000",
    "1101111100110011",
    "1110000000011111",
    "1110000101100010",
    "1110001011101111",
    "1110010010100111",
    "1110011001110101",
    "1110100001000101",
    "1110101000010000",
    "1110101111011010",
    "1110110110100101",
    "1110111101110011",
    "1111000101000000",
    "1111001011111101",
    "1111010010011100",
    "1111011000001100",
    "1111011101001010",
    "1111100001010111",
    "1111100100111011",
    "1111101000001000",
    "1111101011001101",
    "1111101110010100",
    "1111110001100001",
    "1111110100110001",
    "1111110111110111",
    "1111111010101000",
    "1111111100110101",
    "1111111110010101",
    "1111111111000011",
    "1111111111000000",
    "1111111110010011",
    "1111111101000100",
    "1111111011001111",
    "1111111000101000",
    "1111110100111100",
    "1111101111110101",
    "1111101001001110",
    "1111100001001111",
    "1111011000010000",
    "1111001110110001",
    "1111000101100000",
    "1110111101001010",
    "1110110110100010",
    "1110110010010000",
    "1110110000110001",
    "1110110010001101",
    "1110110110011000",
    "1110111100101011",
    "1111000100010010",
    "1111001100010110",
    "1111010100001010",
    "1111011011001110",
    "1111100001010101",
    "1111100110011110",
    "1111101010101010",
    "1111101101111101",
    "1111110000010110",
    "1111110001110010",
    "1111110010001011",
    "1111110001011101",
    "1111101111100111",
    "1111101100101101",
    "1111101000111000",
    "1111100100001101",
    "1111011110110001",
    "1111011000101010",
    "1111010001111001",
    "1111001010101010",
    "1111000011001011",
    "1110111100000001",
    "1110110101110110",
    "1110110001010100",
    "1110101110111010",
    "1110101110101101",
    "1110110000011100",
    "1110110011100001",
    "1110110111010101",
    "1110111011011011",
    "1110111111101000",
    "1111000011111100",
    "1111001000101111",
    "1111001110010100",
    "1111010100111011",
    "1111011100101110",
    "1111100101100100",
    "1111101111000010",
    "1111111000011101",
    "1111111110111100",
    "1111110111111111",
    "1111110011000111",
    "1111110000011101",
    "1111101111110011",
    "1111110000101001",
    "1111110010100001",
    "1111110101000000",
    "1111110111111111",
    "1111111011100011",
    "1111111111110111",
    "1111111010110110",
    "1111110100100111",
    "1111101101100111",
    "1111100110011000",
    "1111011111101000",
    "1111011010000110",
    "1111010110010000",
    "1111010100010011",
    "1111010011111110",
    "1111010100110011",
    "1111010110001110",
    "1111010111111100",
    "1111011001110111",
    "1111011100001100",
    "1111011111000111",
    "1111100010110100",
    "1111100111010110",
    "1111101100100100",
    "1111110010011000",
    "1111111000100110",
    "1111111111000010",
    "1111111010100011",
    "1111110100100100",
    "1111101111011000",
    "1111101011010100",
    "1111101000100100",
    "1111100111001101",
    "1111100111010000",
    "1111101000101111",
    "1111101011101011",
    "1111110000000011",
    "1111110101100111",
    "1111111011110110",
    "1111111110000010",
    "1111111000111100",
    "1111110101100011",
    "1111110100001010",
    "1111110100101010",
    "1111110110100010",
    "1111111001000100",
    "1111111011011101",
    "1111111101000101",
    "1111111101100010",
    "1111111100101010",
    "1111111010100100",
    "1111110111011111",
    "1111110011110000",
    "1111101111110001",
    "1111101011110111",
    "1111101000010010",
    "1111100101010000",
    "1111100010111011",
    "1111100001011110",
    "1111100001000011",
    "1111100001111001",
    "1111100100001011",
    "1111101000000001",
    "1111101101010111",
    "1111110011111101",
    "1111111011011111",
    "1111111100011111",
    "1111110100100000",
    "1111101100111101",
    "1111100110010000",
    "1111100000101011",
    "1111011100100001",
    "1111011001111100",
    "1111011000111110",
    "1111011001010110",
    "1111011010101011",
    "1111011100010110",
    "1111011101101011",
    "1111011110001010",
    "1111011101100110",
    "1111011100001100",
    "1111011010100011",
    "1111011001010101",
    "1111011001000111",
    "1111011010010011",
    "1111011100110010",
    "1111100000001111",
    "1111100100000110",
    "1111100111101100",
    "1111101010011001",
    "1111101011110100",
    "1111101011111001",
    "1111101010110100",
    "1111101000111110",
    "1111100110110111",
    "1111100100111011",
    "1111100011011000",
    "1111100010010111",
    "1111100001110110",
    "1111100001101100",
    "1111100001110001",
    "1111100001111101",
    "1111100010000010",
    "1111100001110000",
    "1111100000111000",
    "1111011111001100",
    "1111011100011011",
    "1111011000011101",
    "1111010011000011",
    "1111001011111101",
    "1111000011001111",
    "1110111001001011",
    "1110101110100001",
    "1110100100010011",
    "1110011011100101",
    "1110010101000101",
    "1110010001000000",
    "1110001110111101",
    "1110001110000111",
    "1110001101101011",
    "1110001101000111",
    "1110001100010110",
    "1110001011101010",
    "1110001011100000",
    "1110001100011001",
    "1110001110101011",
    "1110010010011101",
    "1110010111101010",
    "1110011101111010",
    "1110100100101001",
    "1110101011001001",
    "1110110000101011",
    "1110110100100111",
    "1110110110101000",
    "1110110110110100",
    "1110110101100101",
    "1110110011101001",
    "1110110001110001",
    "1110110000100110",
    "1110110000100011",
    "1110110001110110",
    "1110110100100100",
    "1110111000110000",
    "1110111110011111",
    "1111000101110110",
    "1111001110110110",
    "1111011001100010",
    "1111100101100101",
    "1111110010100011",
    "1111111111101011",
    "1111110011111000",
    "1111101000111100",
    "1111100000000010",
    "1111011001010011",
    "1111010100100010",
    "1111010001010000",
    "1111001111000100",
    "1111001101100110",
    "1111001100101101",
    "1111001100011011",
    "1111001100110111",
    "1111001110000000",
    "1111001111110011",
    "1111010010000110",
    "1111010100101100",
    "1111010111011111",
    "1111011010010011",
    "1111011101000101",
    "1111011111110000",
    "1111100010001000",
    "1111100100000110",
    "1111100101100101",
    "1111100110101001",
    "1111100111011010",
    "1111101000000011",
    "1111101000110001",
    "1111101001101100",
    "1111101010110110",
    "1111101100001010",
    "1111101101100011",
    "1111101110111100",
    "1111110000001111",
    "1111110001010100",
    "1111110010000110",
    "1111110010011011",
    "1111110010010001",
    "1111110001101000",
    "1111110000100100",
    "1111101111010011",
    "1111101110001001",
    "1111101101010111",
    "1111101101001001",
    "1111101101100100",
    "1111101110011100",
    "1111101111011111",
    "1111110000010100",
    "1111110000101111",
    "1111110000101001",
    "1111110000010011",
    "1111110000000100",
    "1111110000011010",
    "1111110001110010",
    "1111110100011101",
    "1111111000011011",
    "1111111101101001",
    "1111111100000100",
    "1111110100111000",
    "1111101100110100",
    "1111100011111011",
    "1111011010011101",
    "1111010000110000",
    "1111000111011011",
    "1110111111000100",
    "1110111000001001",
    "1110110010111001",
    "1110101111001111",
    "1110101100110010",
    "1110101011000110",
    "1110101001110101",
    "1110101000111010",
    "1110101000011010",
    "1110101000011110",
    "1110101001010110",
    "1110101011000100",
    "1110101101100000",
    "1110110000011110",
    "1110110011101001",
    "1110110110110001",
    "1110111001101000",
    "1110111100001001",
    "1110111110010001",
    "1111000000000000",
    "1111000001011010",
    "1111000010100001",
    "1111000011010111",
    "1111000011111001",
    "1111000100001010",
    "1111000100001010",
    "1111000011111001",
    "1111000011011000",
    "1111000010100100",
    "1111000001011100",
    "1111000000000000",
    "1110111110010001",
    "1110111100010110",
    "1110111010011001",
    "1110111000101101",
    "1110110111100111",
    "1110110111011011",
    "1110111000010110",
    "1110111010100000",
    "1110111101110111",
    "1111000010010000",
    "1111000111100000",
    "1111001101100011",
    "1111010100010011",
    "1111011011110101",
    "1111100100001010",
    "1111101101010001",
    "1111110111001010",
    "1111111110010100",
    "1111110011010100",
    "1111100111111110",
    "1111011100100001",
    "1111010001011111",
    "1111000111100000",
    "1110111111010100",
    "1110111001101010",
    "1110110110111110",
    "1110110111011010",
    "1110111010110000",
    "1111000000011110",
    "1111000111101100",
    "1111001111011100",
    "1111010110101101",
    "1111011100100110",
    "1111100000010111",
    "1111100001100100",
    "1111100000001100",
    "1111011100100001",
    "1111010111001011",
    "1111010000111001",
    "1111001010011011",
    "1111000100011000",
    "1110111111001010",
    "1110111010111101",
    "1110110111101111",
    "1110110101011010",
    "1110110011110011",
    "1110110010101110",
    "1110110001111001",
    "1110110000111101",
    "1110101111010111",
    "1110101100110000",
    "1110101000111111",
    "1110100100010010",
    "1110011111000111",
    "1110011010001100",
    "1110010110010101",
    "1110010100000101",
    "1110010011101110",
    "1110010101011000",
    "1110011000111001",
    "1110011110000101",
    "1110100100101010",
    "1110101100011001",
    "1110110100110111",
    "1110111101101000",
    "1111000110000110",
    "1111001101110010",
    "1111010100010010",
    "1111011001011000",
    "1111011101000100",
    "1111011111011001",
    "1111100000100001",
    "1111100000011111",
    "1111011111010110",
    "1111011101000101",
    "1111011001110100",
    "1111010101100100",
    "1111010000100001",
    "1111001010111000",
    "1111000100111100",
    "1110111111000010",
    "1110111001011101",
    "1110110100100100",
    "1110110000100011",
    "1110101101100001",
    "1110101011100000",
    "1110101010011000",
    "1110101010001001",
    "1110101010110010",
    "1110101100010110",
    "1110101110111011",
    "1110110010011111",
    "1110110110111100",
    "1110111100000010",
    "1111000001011111",
    "1111000111000001",
    "1111001100010111",
    "1111010001011110",
    "1111010110010000",
    "1111011010110111",
    "1111011111010111",
    "1111100011101111",
    "1111100111110111",
    "1111101011010111",
    "1111101101110000",
    "1111101110100100",
    "1111101101011001",
    "1111101010001000",
    "1111100101000001",
    "1111011110101011",
    "1111010111110100",
    "1111010001001111",
    "1111001011100011",
    "1111000111000011",
    "1111000011101111",
    "1111000001011110",
    "1110111111111101",
    "1110111111000000",
    "1110111110100110",
    "1110111110110110",
    "1111000000000010",
    "1111000010010101",
    "1111000101111001",
    "1111001010101111",
    "1111010000101100",
    "1111010111011011",
    "1111011110011001",
    "1111100100110111",
    "1111101010001100",
    "1111101101110000",
    "1111101111010000",
    "1111101110110001",
    "1111101100110010",
    "1111101010001000",
    "1111100111110011",
    "1111100110101010",
    "1111100111011000",
    "1111101010001111",
    "1111101111000010",
    "1111110101010000",
    "1111111100000111",
    "1111111101001000",
    "1111110111001111",
    "1111110010100100",
    "1111101111001111",
    "1111101101000111",
    "1111101100000011",
    "1111101011111011",
    "1111101100110011",
    "1111101110110110",
    "1111110010010011",
    "1111110111010110",
    "1111111101111001",
    "1111111010001110",
    "1111110001100000",
    "1111101000100000",
    "1111011111110000",
    "1111010111110010",
    "1111010000111110",
    "1111001011101000",
    "1111000111101111",
    "1111000101010000",
    "1111000011111100",
    "1111000011101100",
    "1111000100011000",
    "1111000110000011",
    "1111001000111001",
    "1111001101000111",
    "1111010010111001",
    "1111011010011011",
    "1111100011101001",
    "1111101110010100",
    "1111111001111111",
    "1111111001111100",
    "1111101110011000",
    "1111100100000110",
    "1111011011110010",
    "1111010110000000",
    "1111010010111011",
    "1111010010011111",
    "1111010100010010",
    "1111010111101010",
    "1111011011111010",
    "1111100000010111",
    "1111100100011100",
    "1111100111101100",
    "1111101001111000",
    "1111101010110010",
    "1111101010010111",
    "1111101000101100",
    "1111100101111110",
    "1111100010101001",
    "1111011111001101",
    "1111011100001110",
    "1111011010000100",
    "1111011000111110",
    "1111011000111001",
    "1111011001101010",
    "1111011010111100",
    "1111011100010110",
    "1111011101100001",
    "1111011110001100",
    "1111011110001010",
    "1111011101011100",
    "1111011100000111",
    "1111011010011000",
    "1111011000011010",
    "1111010110010011",
    "1111010100000011",
    "1111010001011100",
    "1111001110010100",
    "1111001010011110",
    "1111000101111011",
    "1111000000111001",
    "1110111011110101",
    "1110110111010001",
    "1110110011110110",
    "1110110010000011",
    "1110110010010000",
    "1110110100100100",
    "1110111000110010",
    "1110111110100011",
    "1111000101011000",
    "1111001100110011",
    "1111010100011111",
    "1111011100000100",
    "1111100011010000",
    "1111101001110001",
    "1111101111010011",
    "1111110011100111",
    "1111110110100100",
    "1111111000001001",
    "1111111000100001",
    "1111110111111000",
    "1111110110011100",
    "1111110100010001",
    "1111110001011101",
    "1111101110000010",
    "1111101010001011",
    "1111100110001000",
    "1111100010001000",
    "1111011110011001",
    "1111011010111000",
    "1111010111010101",
    "1111010011010010",
    "1111001110001001",
    "1111000111011000",
    "1110111110101011",
    "1110110011111000",
    "1110100111010011",
    "1110011001100010",
    "1110001011100101",
    "1101111110100011",
    "1101110011100111",
    "1101101011100000",
    "1101100110101000",
    "1101100100111100",
    "1101100110001001",
    "1101101001110100",
    "1101101111100011",
    "1101110111000110",
    "1110000000010101",
    "1110001011000111",
    "1110010111000110",
    "1110100011111001",
    "1110110000111101",
    "1110111101101101",
    "1111001001101010",
    "1111010100011010",
    "1111011101110000",
    "1111100101100010",
    "1111101011110000",
    "1111110000100000",
    "1111110011111010",
    "1111110110001100",
    "1111110111101000",
    "1111111000011011",
    "1111111000101110",
    "1111111000101001",
    "1111111000010000",
    "1111110111101011",
    "1111110111000101",
    "1111110110101011",
    "1111110110101011",
    "1111110111001011",
    "1111111000001010",
    "1111111001100010",
    "1111111011000101",
    "1111111100100011",
    "1111111101110101",
    "1111111110111000",
    "1111111111110111",
    "1111111110111010",
    "1111111101001000",
    "1111111010011111",
    "1111110110110000",
    "1111110001111010",
    "1111101100001101",
    "1111100110000110",
    "1111100000001000",
    "1111011010110101",
    "1111010110100000",
    "1111010011010000",
    "1111010000110011",
    "1111001110110001",
    "1111001100110010",
    "1111001010100011",
    "1111000111111111",
    "1111000101010011",
    "1111000010101110",
    "1111000000100111",
    "1110111111010010",
    "1110111110110110",
    "1110111111011001",
    "1111000000110011",
    "1111000010111011",
    "1111000101100111",
    "1111001000101000",
    "1111001011110000",
    "1111001110110000",
    "1111010001100001",
    "1111010011111011",
    "1111010101111110",
    "1111010111101111",
    "1111011001011000",
    "1111011011000010",
    "1111011100110000",
    "1111011110011111",
    "1111100000000010",
    "1111100001000101",
    "1111100001010100",
    "1111100000100100",
    "1111011110111101",
    "1111011100101110",
    "1111011010011000",
    "1111011000100010",
    "1111010111101010",
    "1111011000001001",
    "1111011010001011",
    "1111011101101000",
    "1111100010011100",
    "1111101000010111",
    "1111101111011000",
    "1111110111100000",
    "1111111111001011",
    "1111110100110110",
    "1111101001110001",
    "1111011110011110",
    "1111010011100100",
    "1111001001100101",
    "1111000000110000",
    "1110111001000010",
    "1110110010001111",
    "1110101100000010",
    "1110100110010101",
    "1110100001001000",
    "1110011100101000",
    "1110011001000111",
    "1110010110101101",
    "1110010101011111",
    "1110010101010111",
    "1110010110001110",
    "1110010111111110",
    "1110011010100011",
    "1110011101111101",
    "1110100001111110",
    "1110100110010101",
    "1110101010100101",
    "1110101110010010",
    "1110110001010000",
    "1110110011100001",
    "1110110101010010",
    "1110110110111110",
    "1110111000111100",
    "1110111011011001",
    "1110111110010111",
    "1111000001101011",
    "1111000101000001",
    "1111001000001000",
    "1111001010101111",
    "1111001100110010",
    "1111001110010110",
    "1111001111101000",
    "1111010000111001",
    "1111010010100110",
    "1111010100111011",
    "1111011000000100",
    "1111011011111000",
    "1111100000000011",
    "1111100011111110",
    "1111100111000011",
    "1111101000101110",
    "1111101000101100",
    "1111100111000100",
    "1111100100010000",
    "1111100000111011",
    "1111011101110011",
    "1111011011100101",
    "1111011010101111",
    "1111011011100001",
    "1111011110000100",
    "1111100010010101",
    "1111101000010100",
    "1111110000000001",
    "1111111001011010",
    "1111111011100001",
    "1111101110111011",
    "1111100001000000",
    "1111010010001010",
    "1111000010111110",
    "1110110100010011",
    "1110100110111110",
    "1110011011101101",
    "1110010010111101",
    "1110001100110101",
    "1110001001000110",
    "1110000111010110",
    "1110000111001001",
    "1110001000000001",
    "1110001001101010",
    "1110001011110000",
    "1110001101111101",
    "1110010000000000",
    "1110010001101011",
    "1110010010110011",
    "1110010011010011",
    "1110010011010111",
    "1110010011001011",
    "1110010011001101",
    "1110010011111011",
    "1110010101111110",
    "1110011001111101",
    "1110100000011100",
    "1110101001101010",
    "1110110101011111",
    "1111000011010111",
    "1111010010001000",
    "1111100000010111",
    "1111101100100100",
    "1111110101101110",
    "1111111011011101",
    "1111111110001010",
    "1111111110101010",
    "1111111110000011",
    "1111111101001011",
    "1111111100100001",
    "1111111100000110",
    "1111111011101101",
    "1111111011000111",
    "1111111010001110",
    "1111111001000111",
    "1111110111111000",
    "1111110110100000",
    "1111110100110101",
    "1111110010100110",
    "1111101111101001",
    "1111101100000001",
    "1111101000001001",
    "1111100100100111",
    "1111100001111101",
    "1111100000010111",
    "1111011111101011",
    "1111011111011001",
    "1111011110111010",
    "1111011101110011",
    "1111011100000010",
    "1111011001111100",
    "1111011000001001",
    "1111010111010000",
    "1111010111101101",
    "1111011001101101",
    "1111011101001100",
    "1111100001110110",
    "1111100111001101",
    "1111101100101110",
    "1111110001110001",
    "1111110101101011",
    "1111110111111000",
    "1111110111111101",
    "1111110101101111",
    "1111110001010101",
    "1111101011000000",
    "1111100011000110",
    "1111011001111101",
    "1111001111111111",
    "1111000101100100",
    "1110111011010001",
    "1110110001111000",
    "1110101010000111",
    "1110100100100100",
    "1110100001011111",
    "1110100000111000",
    "1110100010010111",
    "1110100101011101",
    "1110101001101011",
    "1110101110110000",
    "1110110100100100",
    "1110111011000111",
    "1111000010011010",
    "1111001010011000",
    "1111010010111001",
    "1111011011101101",
    "1111100100100000",
    "1111101100111010",
    "1111110100100000",
    "1111111010111111",
    "1111111111110110",
    "1111111100001010",
    "1111111001110010",
    "1111111000100000",
    "1111111000000001",
    "1111111000000111",
    "1111111000101001",
    "1111111001101100",
    "1111111011011110",
    "1111111110010110",
    "1111111101010001",
    "1111110111001011",
    "1111101111010101",
    "1111100110000110",
    "1111011100010001",
    "1111010010111110",
    "1111001011010100",
    "1111000110001000",
    "1111000011110011",
    "1111000100000110",
    "1111000110011010",
    "1111001001111010",
    "1111001101110010",
    "1111010001010010",
    "1111010100000001",
    "1111010101110111",
    "1111010110110111",
    "1111010111010000",
    "1111010111011010",
    "1111010111110111",
    "1111011001000111",
    "1111011011100001",
    "1111011111010010",
    "1111100100010101",
    "1111101010011010",
    "1111110001000101",
    "1111110111111100",
    "1111111110100011",
    "1111111011010111",
    "1111110110001100",
    "1111110010001000",
    "1111101111011010",
    "1111101110001100",
    "1111101110100100",
    "1111110000100000",
    "1111110011110111",
    "1111111000010101",
    "1111111101100010",
    "1111111100111111",
    "1111110111110001",
    "1111110011000011",
    "1111101111000001",
    "1111101011100011",
    "1111101000011100",
    "1111100101011111",
    "1111100010100001",
    "1111011111011111",
    "1111011100101000",
    "1111011010001100",
    "1111011000100010",
    "1111010111111010",
    "1111011000100011",
    "1111011010011011",
    "1111011101011100",
    "1111100001011010",
    "1111100110001001",
    "1111101011011101",
    "1111110001000011",
    "1111110110110000",
    "1111111100010100",
    "1111111110011010",
    "1111111001100110",
    "1111110101000110",
    "1111110000110001",
    "1111101100011010",
    "1111100111110101",
    "1111100011000101",
    "1111011110010010",
    "1111011001110111",
    "1111010110001011",
    "1111010011100110",
    "1111010010010101",
    "1111010010100001",
    "1111010011111100",
    "1111010110011111",
    "1111011001110010",
    "1111011101100110",
    "1111100001101100",
    "1111100101110111",
    "1111101001111000",
    "1111101101011001",
    "1111110000001000",
    "1111110001110100",
    "1111110010010010",
    "1111110001100100",
    "1111101111110111",
    "1111101101100001",
    "1111101010111001",
    "1111101000010100",
    "1111100101111100",
    "1111100011111001",
    "1111100010001011",
    "1111100000110101",
    "1111011111110110",
    "1111011111010010",
    "1111011111001000",
    "1111011111010111",
    "1111011111110101",
    "1111100000001111",
    "1111100000010010",
    "1111011111100110",
    "1111011101110111",
    "1111011010101101",
    "1111010101110111",
    "1111001111000111",
    "1111000110010010",
    "1110111011100001",
    "1110101111011001",
    "1110100010101111",
    "1110010110110010",
    "1110001100101011",
    "1110000101001110",
    "1110000000110101",
    "1101111111001111",
    "1101111111111010",
    "1110000010000110",
    "1110000101001110",
    "1110001000111010",
    "1110001100111111",
    "1110010001010100",
    "1110010101101100",
    "1110011001110101",
    "1110011101010110",
    "1110011111110011",
    "1110100000111110",
    "1110100000110000",
    "1110011111001111",
    "1110011100101011",
    "1110011001011101",
    "1110010101111110",
    "1110010010110001",
    "1110010000011100",
    "1110001111100011",
    "1110010000100011",
    "1110010011101100",
    "1110011001000100",
    "1110100000100011",
    "1110101001111010",
    "1110110100110111",
    "1111000001000011",
    "1111001110000000",
    "1111011011001010",
    "1111100111110110",
    "1111110011011000",
    "1111111101001110",
    "1111111010110110",
    "1111110100110100",
    "1111110000010011",
    "1111101100110100",
    "1111101001110100",
    "1111100111000000",
    "1111100100001110",
    "1111100001100111",
    "1111011111011001",
    "1111011101101011",
    "1111011100101010",
    "1111011100010001",
    "1111011100011110",
    "1111011101001100",
    "1111011110010100",
    "1111011111110011",
    "1111100001101001",
    "1111100011110011",
    "1111100110001101",
    "1111101000110001",
    "1111101011011010",
    "1111101110000000",
    "1111110000011010",
    "1111110010100000",
    "1111110100001010",
    "1111110101010001",
    "1111110101110111",
    "1111110110000000",
    "1111110101111000",
    "1111110101101100",
    "1111110101100111",
    "1111110101110000",
    "1111110110001000",
    "1111110110101000",
    "1111110111001100",
    "1111110111101100",
    "1111111000000001",
    "1111111000000011",
    "1111110111101011",
    "1111110110110010",
    "1111110101011011",
    "1111110011101000",
    "1111110001100111",
    "1111101111100010",
    "1111101101100100",
    "1111101011110100",
    "1111101010010000",
    "1111101000111001",
    "1111100111101110",
    "1111100110110100",
    "1111100110010011",
    "1111100110011101",
    "1111100111011111",
    "1111101001101100",
    "1111101101010011",
    "1111110010100110",
    "1111111001110001",
    "1111111101000101",
    "1111110010001001",
    "1111100101110111",
    "1111011001000110",
    "1111001100111000",
    "1111000010001101",
    "1110111001111010",
    "1110110100010101",
    "1110110001011001",
    "1110110000011111",
    "1110110000111101",
    "1110110010000110",
    "1110110011011010",
    "1110110100100111",
    "1110110101101100",
    "1110110110101000",
    "1110110111100101",
    "1110111000100010",
    "1110111001100000",
    "1110111010100000",
    "1110111011100110",
    "1110111100111010",
    "1110111110101001",
    "1111000000111110",
    "1111000011111000",
    "1111000111001101",
    "1111001010100010",
    "1111001101011011",
    "1111001111010100",
    "1111001111111010",
    "1111001110111111",
    "1111001100101011",
    "1111001001011001",
    "1111000101101010",
    "1111000001111110",
    "1110111110110011",
    "1110111100011110",
    "1110111011000010",
    "1110111010011001",
    "1110111010010110",
    "1110111010110000",
    "1110111011100001",
    "1110111100110111",
    "1110111110111111",
    "1111000010010000",
    "1111000111000001",
    "1111001101010010",
    "1111010100111011",
    "1111011101011100",
    "1111100110010011",
    "1111101110111010",
    "1111110110101111",
    "1111111101100011",
    "1111111100100110",
    "1111110111011111",
    "1111110010101100",
    "1111101101101100",
    "1111101000001011",
    "1111100010000011",
    "1111011011100011",
    "1111010101001001",
    "1111001111011001",
    "1111001010110000",
    "1111000111100011",
    "1111000101110100",
    "1111000101011000",
    "1111000110001000",
    "1111000111110101",
    "1111001010011011",
    "1111001101101000",
    "1111010001001010",
    "1111010100011111",
    "1111010111000001",
    "1111011000001011",
    "1111010111101100",
    "1111010101011111",
    "1111010001110011",
    "1111001101000000",
    "1111000111100011",
    "1111000001101110",
    "1110111011101101",
    "1110110101101110",
    "1110101111110101",
    "1110101010010001",
    "1110100101001101",
    "1110100000110110",
    "1110011101010111",
    "1110011010110111",
    "1110011001011000",
    "1110011000110101",
    "1110011001010000",
    "1110011010011110",
    "1110011100010111",
    "1110011110111010",
    "1110100010000000",
    "1110100101101110",
    "1110101010000001",
    "1110101110111000",
    "1110110100001101",
    "1110111001101111",
    "1110111111001010",
    "1111000100001010",
    "1111001000011101",
    "1111001100000001",
    "1111001110110101",
    "1111010001000011",
    "1111010010111000",
    "1111010100011101",
    "1111010101110110",
    "1111010111000001",
    "1111010111110101",
    "1111010111111111",
    "1111010111010000",
    "1111010101010011",
    "1111010010000000",
    "1111001101010110",
    "1111000111011111",
    "1111000000101100",
    "1110111001011011",
    "1110110010001010",
    "1110101011011101",
    "1110100101101111",
    "1110100001011110",
    "1110011110111111",
    "1110011110100100",
    "1110100000011010",
    "1110100100100100",
    "1110101010111000",
    "1110110010111110",
    "1110111100010011",
    "1111000110000011",
    "1111001111011001",
    "1111010111100111",
    "1111011110001100",
    "1111100010111110",
    "1111100110000011",
    "1111100111110011",
    "1111101000101111",
    "1111101001010000",
    "1111101001101001",
    "1111101001111100",
    "1111101001111100",
    "1111101001010111",
    "1111100111111101",
    "1111100101100010",
    "1111100010001010",
    "1111011101111111",
    "1111011001010101",
    "1111010100100000",
    "1111001111110110",
    "1111001011100101",
    "1111000111111110",
    "1111000101001000",
    "1111000011001010",
    "1111000010000011",
    "1111000001110100",
    "1111000010011010",
    "1111000011111000",
    "1111000110001110",
    "1111001001100011",
    "1111001101110011",
    "1111010010101111",
    "1111010111110111",
    "1111011100101000",
    "1111100000011010",
    "1111100010110100",
    "1111100011100111",
    "1111100010111110",
    "1111100001010100",
    "1111011111010111",
    "1111011101111011",
    "1111011101110111",
    "1111011111101110",
    "1111100011110110",
    "1111101010001000",
    "1111110010001001",
    "1111111011001010",
    "1111111011100100",
    "1111110010110101",
    "1111101011000111",
    "1111100100101100",
    "1111011111101100",
    "1111011100000111",
    "1111011001111010",
    "1111011001000111",
    "1111011001110111",
    "1111011100001111",
    "1111100000011010",
    "1111100110011101",
    "1111101110011000",
    "1111111000001000",
    "1111111100011110",
    "1111110000000101",
    "1111100011100001",
    "1111010111110111",
    "1111001110001100",
    "1111000111010101",
    "1111000011101010",
    "1111000011000110",
    "1111000101000110",
    "1111001000111100",
    "1111001101111101",
    "1111010011100111",
    "1111011001101011",
    "1111100000000101",
    "1111100110110101",
    "1111101101110111",
    "1111110101000000",
    "1111111011111000",
    "1111111101110111",
    "1111111000101111",
    "1111110101000010",
    "1111110010111111",
    "1111110010101001",
    "1111110011111001",
    "1111110110011100",
    "1111111001110010",
    "1111111101010011",
    "1111111111101000",
    "1111111101101000",
    "1111111100111101",
    "1111111101110001",
    "1111111111111111",
    "1111111100100011",
    "1111111000000110",
    "1111110010110011",
    "1111101100110111",
    "1111100110101000",
    "1111100000100100",
    "1111011011010011",
    "1111010111011010",
    "1111010101010111",
    "1111010101001110",
    "1111010110101100",
    "1111011001000010",
    "1111011011011101",
    "1111011101000100",
    "1111011101010001",
    "1111011011111000",
    "1111011000111110",
    "1111010100111001",
    "1111010000001100",
    "1111001011011110",
    "1111000111001110",
    "1111000011110100",
    "1111000001011100",
    "1110111111111101",
    "1110111111001100",
    "1110111110110011",
    "1110111110011111",
    "1110111110001001",
    "1110111101110010",
    "1110111101101110",
    "1110111110011100",
    "1111000000010100",
    "1111000011101001",
    "1111001000010110",
    "1111001110001111",
    "1111010100110110",
    "1111011011101010",
    "1111100010010101",
    "1111101000101010",
    "1111101110100100",
    "1111110100000010",
    "1111111001000101",
    "1111111101101101",
    "1111111110001001",
    "1111111010101010",
    "1111110111111011",
    "1111110110000001",
    "1111110101000001",
    "1111110100111101",
    "1111110101110011",
    "1111110111100101",
    "1111111010011010",
    "1111111110010110",
    "1111111100011011",
    "1111110101111010",
    "1111101110000100",
    "1111100100111001",
    "1111011010100101",
    "1111001111010110",
    "1111000011100001",
    "1110110111100011",
    "1110101011111101",
    "1110100001001111",
    "1110010111110010",
    "1110001111110110",
    "1110001001011101",
    "1110000100011010",
    "1110000000100011",
    "1101111101101000",
    "1101111011101000",
    "1101111010100110",
    "1101111010110100",
    "1101111100011110",
    "1101111111110000",
    "1110000100101100",
    "1110001011001010",
    "1110010010111101",
    "1110011011101111",
    "1110100101001110",
    "1110101111000111",
    "1110111001000110",
    "1111000010110011",
    "1111001011110111",
    "1111010011111011",
    "1111011010101011",
    "1111100000000111",
    "1111100100001011",
    "1111100111001001",
    "1111101001001110",
    "1111101010101110",
    "1111101011111000",
    "1111101100110110",
    "1111101101110010",
    "1111101110110000",
    "1111101111110100",
    "1111110001000000",
    "1111110010010101",
    "1111110011110010",
    "1111110101010100",
    "1111110110110101",
    "1111111000001100",
    "1111111001010100",
    "1111111010000101",
    "1111111010100001",
    "1111111010110001",
    "1111111011000100",
    "1111111011110000",
    "1111111101001000",
    "1111111111011001",
    "1111111101011011",
    "1111111001100110",
    "1111110101010100",
    "1111110000111001",
    "1111101100011100",
    "1111100111111101",
    "1111100011010111",
    "1111011110100110",
    "1111011001101000",
    "1111010100100000",
    "1111001111011010",
    "1111001010100101",
    "1111000110001110",
    "1111000010100111",
    "1111000000000010",
    "1110111110101000",
    "1110111110011111",
    "1110111111101100",
    "1111000010000110",
    "1111000101011011",
    "1111001001010101",
    "1111001101010110",
    "1111010001001101",
    "1111010100101010",
    "1111010111101000",
    "1111011010001100",
    "1111011100011011",
    "1111011110011110",
    "1111100000010101",
    "1111100001111110",
    "1111100011010000",
    "1111100011111100",
    "1111100011111100",
    "1111100011001101",
    "1111100001110011",
    "1111011111111011",
    "1111011101111010",
    "1111011100000001",
    "1111011010100011",
    "1111011001101111",
    "1111011001101010",
    "1111011010011011",
    "1111011100000100",
    "1111011110100011",
    "1111100001110001",
    "1111100101101001",
    "1111101010000100",
    "1111101111000101",
    "1111110100111001",
    "1111111011101110",
    "1111111100001100",
    "1111110010110110",
    "1111101000011011",
    "1111011101011001",
    "1111010010010100",
    "1111000111101010",
    "1110111101111000",
    "1110110101000110",
    "1110101101011011",
    "1110100110110100",
    "1110100001011001",
    "1110011101010001",
    "1110011010100101",
    "1110011001011110",
    "1110011001111010",
    "1110011011101111",
    "1110011110101000",
    "1110100010001010",
    "1110100101111001",
    "1110101001010110",
    "1110101100001001",
    "1110101101111111",
    "1110101110110000",
    "1110101110011111",
    "1110101101011011",
    "1110101011111010",
    "1110101010011011",
    "1110101001100000",
    "1110101001100010",
    "1110101010101010",
    "1110101100110011",
    "1110101111110000",
    "1110110011000110",
    "1110110110100010",
    "1110111001111100",
    "1110111101010110",
    "1111000000110110",
    "1111000100100111",
    "1111001000100011",
    "1111001100011100",
    "1111001111111111",
    "1111010010101111",
    "1111010100100000",
    "1111010101001101",
    "1111010100111001",
    "1111010011110110",
    "1111010010010111",
    "1111010000101100",
    "1111001111001000",
    "1111001101111000",
    "1111001101001010",
    "1111001101001111",
    "1111001110011001",
    "1111010000110101",
    "1111010100101010",
    "1111011001111101",
    "1111100000101100",
    "1111101000110101",
    "1111110010010000",
    "1111111100111011",
    "1111110111010111",
    "1111101011000001",
    "1111011110100011",
    "1111010010100001",
    "1111000111011010",
    "1110111101100110",
    "1110110101001001",
    "1110101110000000",
    "1110100111111001",
    "1110100010100010",
    "1110011101101110",
    "1110011001011001",
    "1110010101100000",
    "1110010010001000",
    "1110001111010100",
    "1110001101000101",
    "1110001011100000",
    "1110001010100011",
    "1110001010001111",
    "1110001010100011",
    "1110001011011011",
    "1110001100111010",
    "1110001111000000",
    "1110010001110001",
    "1110010101011000",
    "1110011010000100",
    "1110100000001000",
    "1110100111110111",
    "1110110001010100",
    "1110111100010111",
    "1111001000011011",
    "1111010100100100",
    "1111011111101000",
    "1111101000100011",
    "1111101110101111",
    "1111110010001000",
    "1111110011010011",
    "1111110011000011",
    "1111110010011000",
    "1111110001111000",
    "1111110001110100",
    "1111110010001001",
    "1111110010100001",
    "1111110010100110",
    "1111110010000110",
    "1111110000101111",
    "1111101110010110",
    "1111101010110111",
    "1111100110010110",
    "1111100001000101",
    "1111011011100000",
    "1111010110010010",
    "1111010010000010",
    "1111001111010110",
    "1111001110011111",
    "1111001111011110",
    "1111010001111110",
    "1111010101011111",
    "1111011001010110",
    "1111011101000101",
    "1111100000010001",
    "1111100010101100",
    "1111100100011010",
    "1111100101100111",
    "1111100110101000",
    "1111100111110101",
    "1111101001011110",
    "1111101011100110",
    "1111101110000111",
    "1111110000101011",
    "1111110010110100",
    "1111110100000001",
    "1111110011110010",
    "1111110001110010",
    "1111101101110110",
    "1111100111111000",
    "1111011111111111",
    "1111010110010101",
    "1111001011010011",
    "1110111111100011",
    "1110110011111011",
    "1110101001011110",
    "1110100001000111",
    "1110011011011110",
    "1110011000110000",
    "1110011000101100",
    "1110011010100110",
    "1110011101110011",
    "1110100001110001",
    "1110100110010011",
    "1110101011011110",
    "1110110001101001",
    "1110111001000100",
    "1111000001111001",
    "1111001011111010",
    "1111010110100111",
    "1111100001010000",
    "1111101011000110",
    "1111110011011100",
    "1111111001110110",
    "1111111110001011",
    "1111111111011011",
    "1111111110101011",
    "1111111111000101",
    "1111111111110011",
    "1111111110100000",
    "1111111101001111",
    "1111111100000111",
    "1111111011000001",
    "1111111001101011",
    "1111110111110000",
    "1111110101000000",
    "1111110001010100",
    "1111101100110100",
    "1111100111110011",
    "1111100010100111",
    "1111011101101001",
    "1111011001001100",
    "1111010101011011",
    "1111010010010111",
    "1111010000000000",
    "1111001110001100",
    "1111001100110101",
    "1111001011101111",
    "1111001010110100",
    "1111001010000100",
    "1111001001100101",
    "1111001001100011",
    "1111001010001111",
    "1111001011111010",
    "1111001110110000",
    "1111010010111001",
    "1111011000010011",
    "1111011110111000",
    "1111100110011000",
    "1111101110100011",
    "1111110111000001",
    "1111111111010110",
    "1111111000111000",
    "1111110010001010",
    "1111101100110100",
    "1111101001000011",
    "1111100110111100",
    "1111100110100001",
    "1111100111101110",
    "1111101010100000",
    "1111101110110001",
    "1111110100010111",
    "1111111010111101",
    "1111111101111010",
    "1111110110111000",
    "1111110000011101",
    "1111101011000010",
    "1111100110110100",
    "1111100011101110",
    "1111100001100001",
    "1111011111110101",
    "1111011110010100",
    "1111011100110111",
    "1111011011011110",
    "1111011010010100",
    "1111011001101101",
    "1111011001111010",
    "1111011011001001",
    "1111011101011100",
    "1111100000110000",
    "1111100100111011",
    "1111101001110011",
    "1111101111001100",
    "1111110100111101",
    "1111111010111101",
    "1111111110111010",
    "1111111000110111",
    "1111110010111111",
    "1111101101011011",
    "1111101000010001",
    "1111100011100111",
    "1111011111101000",
    "1111011100100001",
    "1111011010100011",
    "1111011001111101",
    "1111011010110101",
    "1111011101000100",
    "1111100000001111",
    "1111100011110110",
    "1111100111010101",
    "1111101010001101",
    "1111101100001100",
    "1111101101001100",
    "1111101101010010",
    "1111101100101001",
    "1111101011011111",
    "1111101010000100",
    "1111101000100110",
    "1111100111010101",
    "1111100110011000",
    "1111100101110100",
    "1111100101100111",
    "1111100101101001",
    "1111100101101111",
    "1111100101101110",
    "1111100101100010",
    "1111100101001000",
    "1111100100100010",
    "1111100011101111",
    "1111100010101111",
    "1111100001011100",
    "1111011111110000",
    "1111011101100100",
    "1111011010110101",
    "1111010111011011",
    "1111010011010101",
    "1111001110011001",
    "1111001000100011",
    "1111000001110011",
    "1110111010001011",
    "1110110001111001",
    "1110101001100010",
    "1110100001110000",
    "1110011011010100",
    "1110010110110111",
    "1110010100101010",
    "1110010100100111",
    "1110010110001011",
    "1110011000100111",
    "1110011011001111",
    "1110011101100110",
    "1110011111011110",
    "1110100000111011",
    "1110100010000011",
    "1110100011000000",
    "1110100011100111",
    "1110100011101100",
    "1110100010111001",
    "1110100000111110",
    "1110011101110011",
    "1110011001011001",
    "1110010100000110",
    "1110001110010111",
    "1110001000110000",
    "1110000011111011",
    "1110000000011001",
    "1101111110101110",
    "1101111111001100",
    "1110000001111110",
    "1110000111000110",
    "1110001110011111",
    "1110011000000100",
    "1110100011100111",
    "1110110000110101",
    "1110111111001000",
    "1111001101110101",
    "1111011011111101",
    "1111101000100100",
    "1111110010111100",
    "1111111010101111",
    "1111111111110001",
    "1111111100000100",
    "1111111001010001",
    "1111110110101000",
    "1111110011101100",
    "1111110000010111",
    "1111101100111011",
    "1111101001110001",
    "1111100111001100",
    "1111100101010011",
    "1111100100000000",
    "1111100011000001",
    "1111100010000010",
    "1111100000101110",
    "1111011110111010",
    "1111011100100101",
    "1111011001111001",
    "1111010111000011",
    "1111010100011100",
    "1111010010011001",
    "1111010001001111",
    "1111010001001111",
    "1111010010011101",
    "1111010100111100",
    "1111011000100000",
    "1111011100111111",
    "1111100010000101",
    "1111100111100001",
    "1111101100111101",
    "1111110010000101",
    "1111110110100001",
    "1111111010000001",
    "1111111100011010",
    "1111111101101011",
    "1111111101110110",
    "1111111101000110",
    "1111111011100111",
    "1111111001100101",
    "1111110111001011",
    "1111110100100001",
    "1111110001110010",
    "1111101111000011",
    "1111101100011100",
    "1111101010000100",
    "1111100111111110",
    "1111100110001110",
    "1111100100110110",
    "1111100011111000",
    "1111100011001111",
    "1111100010111110",
    "1111100011001000",
    "1111100011110001",
    "1111100101000001",
    "1111100111000100",
    "1111101010000001",
    "1111101110000100",
    "1111110011010100",
    "1111111001111011",
    "1111111101111011",
    "1111110100001001",
    "1111101000101110",
    "1111011100000100",
    "1111001111000100",
    "1111000010111011",
    "1110111000110111",
    "1110110001110110",
    "1110101110010001",
    "1110101101110111",
    "1110101111110110",
    "1110110011010111",
    "1110110111100010",
    "1110111011110101",
    "1111000000000000",
    "1111000011111100",
    "1111000111100101",
    "1111001010110000",
    "1111001101001111",
    "1111001110110110",
    "1111001111011001",
    "1111001110111000",
    "1111001101011100",
    "1111001011011000",
    "1111001000111010",
    "1111000110001110",
    "1111000011011100",
    "1111000000100100",
    "1110111101101101",
    "1110111010111010",
    "1110111000010101",
    "1110110110000110",
    "1110110100010101",
    "1110110011001010",
    "1110110010100110",
    "1110110010100111",
    "1110110011001111",
    "1110110100010010",
    "1110110101101001",
    "1110110111001110",
    "1110111000111010",
    "1110111010110000",
    "1110111100111000",
    "1110111111100110",
    "1111000011001101",
    "1111000111111100",
    "1111001101111101",
    "1111010101001000",
    "1111011101001100",
    "1111100101100111",
    "1111101101111110",
    "1111110101111000",
    "1111111101001011",
    "1111111100000100",
    "1111110101111000",
    "1111110000001100",
    "1111101011000100",
    "1111100110110010",
    "1111100011101001",
    "1111100001111000",
    "1111100001100110",
    "1111100010100111",
    "1111100100100010",
    "1111100110110101",
    "1111101000111111",
    "1111101010100010",
    "1111101011001100",
    "1111101010110011",
    "1111101001010010",
    "1111100110101101",
    "1111100011001000",
    "1111011110101110",
    "1111011001101010",
    "1111010100001110",
    "1111001110101001",
    "1111001001001100",
    "1111000100000101",
    "1110111111010111",
    "1110111011000100",
    "1110110110111111",
    "1110110011000000",
    "1110101110111010",
    "1110101010101101",
    "1110100110100000",
    "1110100010100010",
    "1110011111001000",
    "1110011100100001",
    "1110011010110100",
    "1110011010000111",
    "1110011010011011",
    "1110011011110011",
    "1110011110010001",
    "1110100001110011",
    "1110100110010000",
    "1110101011011001",
    "1110110000110110",
    "1110110110001101",
    "1110111011000111",
    "1110111111011001",
    "1111000011000110",
    "1111000110011000",
    "1111001001100000",
    "1111001100101000",
    "1111001111111000",
    "1111010011001101",
    "1111010110011101",
    "1111011001011011",
    "1111011011111101",
    "1111011101111000",
    "1111011111000101",
    "1111011111100001",
    "1111011111000101",
    "1111011101110000",
    "1111011011011101",
    "1111011000000110",
    "1111010011101010",
    "1111001110001111",
    "1111001000000001",
    "1111000001011111",
    "1110111011001111",
    "1110110110000001",
    "1110110010011101",
    "1110110001000011",
    "1110110001111011",
    "1110110100111100",
    "1110111001101011",
    "1110111111100100",
    "1111000110000000",
    "1111001100011110",
    "1111010010100110",
    "1111011000000100",
    "1111011100101110",
    "1111100000100001",
    "1111100011010101",
    "1111100101001011",
    "1111100101111110",
    "1111100101101010",
    "1111100100001110",
    "1111100001101001",
    "1111011110000000",
    "1111011001100010",
    "1111010100100101",
    "1111001111100100",
    "1111001010111100",
    "1111000111000001",
    "1111000100000011",
    "1111000010001000",
    "1111000001010010",
    "1111000001011100",
    "1111000010100010",
    "1111000100011100",
    "1111000110111111",
    "1111001001111101",
    "1111001101000010",
    "1111001111111010",
    "1111010010010010",
    "1111010100000000",
    "1111010101000000",
    "1111010101010101",
    "1111010101001110",
    "1111010100111001",
    "1111010100011111",
    "1111010100001000",
    "1111010011110100",
    "1111010011011111",
    "1111010011000101",
    "1111010010101111",
    "1111010010101111",
    "1111010011100110",
    "1111010101110100",
    "1111011001111001",
    "1111100000000111",
    "1111101000011001",
    "1111110010010010",
    "1111111101000111",
    "1111111000000111",
    "1111101110011100",
    "1111100110110001",
    "1111100001110011",
    "1111011111111010",
    "1111100001000011",
    "1111100100111011",
    "1111101010111110",
    "1111110010101011",
    "1111111011100001",
    "1111111010110110",
    "1111110000111000",
    "1111100110111011",
    "1111011101011100",
    "1111010100111110",
    "1111001101111011",
    "1111001000100011",
    "1111000100111001",
    "1111000010110011",
    "1111000010000000",
    "1111000010010101",
    "1111000011101010",
    "1111000110000001",
    "1111001001011101",
    "1111001101111011",
    "1111010011010111",
    "1111011001011000",
    "1111011111101001",
    "1111100101101010",
    "1111101010111011",
    "1111101111000111",
    "1111110010000100",
    "1111110011110000",
    "1111110100010111",
    "1111110100001010",
    "1111110011011010",
    "1111110010011100",
    "1111110001011110",
    "1111110000101000",
    "1111110000000010",
    "1111101111101110",
    "1111101111101100",
    "1111101111111111",
    "1111110000100111",
    "1111110001101010",
    "1111110011001010",
    "1111110101001111",
    "1111110111111100",
    "1111111011011001",
    "1111111111101010",
    "1111111011000111",
    "1111110100111110",
    "1111101101111110",
    "1111100110010101",
    "1111011110100011",
    "1111010111010011",
    "1111010001010000",
    "1111001101000100",
    "1111001010111010",
    "1111001010101011",
    "1111001011110111",
    "1111001101101001",
    "1111001111010010",
    "1111010000001000",
    "1111001111111000",
    "1111001110100001",
    "1111001100001110",
    "1111001001010101",
    "1111000110001001",
    "1111000010111011",
    "1110111111110000",
    "1110111100101101",
    "1110111001111001",
    "1110110111100011",
    "1110110110000110",
    "1110110101110010",
    "1110110110111100",
    "1110111001100101",
    "1110111101101000",
    "1111000010110100",
    "1111001000111100",
    "1111001111101100",
    "1111010110111100",
    "1111011110011100",
    "1111100110000000",
    "1111101101011001",
    "1111110100010100",
    "1111111010100000",
    "1111111111101101",
    "1111111100001001",
    "1111111001001111",
    "1111110111100000",
    "1111110110110111",
    "1111110111001010",
    "1111111000010010",
    "1111111010000101",
    "1111111100011101",
    "1111111111010110",
    "1111111101001001",
    "1111111001000100",
    "1111110100010001",
    "1111101110110000",
    "1111101000011110",
    "1111100001100001",
    "1111011001110101",
    "1111010001011110",
    "1111001000010000",
    "1110111110001100",
    "1110110011010000",
    "1110100111110010",
    "1110011100001111",
    "1110010001010100",
    "1110000111100101",
    "1101111111100110",
    "1101111001101000",
    "1101110101101001",
    "1101110011011100",
    "1101110010101111",
    "1101110011010111",
    "1101110101001110",
    "1101111000011010",
    "1101111100111111",
    "1110000011000011",
    "1110001010100000",
    "1110010011001101",
    "1110011100110111",
    "1110100111001000",
    "1110110001100111",
    "1110111011111101",
    "1111000101101111",
    "1111001110011111",
    "1111010101111001",
    "1111011011101000",
    "1111011111101000",
    "1111100001111101",
    "1111100010111110",
    "1111100011000110",
    "1111100010111001",
    "1111100010111001",
    "1111100011100001",
    "1111100100111110",
    "1111100111010011",
    "1111101010010011",
    "1111101101100110",
    "1111110000101101",
    "1111110011000100",
    "1111110100010010",
    "1111110100001001",
    "1111110010101011",
    "1111110000001011",
    "1111101101001011",
    "1111101010010010",
    "1111101000000110",
    "1111100111000100",
    "1111100111011101",
    "1111101001010011",
    "1111101100011101",
    "1111110000101101",
    "1111110101110101",
    "1111111011101000",
    "1111111110000001",
    "1111110111010110",
    "1111110000100011",
    "1111101001111100",
    "1111100011110001",
    "1111011110010001",
    "1111011001100101",
    "1111010101101110",
    "1111010010100010",
    "1111001111111111",
    "1111001101111101",
    "1111001100011110",
    "1111001011101000",
    "1111001011100001",
    "1111001100010011",
    "1111001101111011",
    "1111010000010101",
    "1111010011010000",
    "1111010110011010",
    "1111011001011101",
    "1111011100001100",
    "1111011110011111",
    "1111100000010010",
    "1111100001100010",
    "1111100010010000",
    "1111100010011010",
    "1111100001111110",
    "1111100000111101",
    "1111011111010110",
    "1111011101001110",
    "1111011010101011",
    "1111010111111001",
    "1111010101000011",
    "1111010010011100",
    "1111010000010010",
    "1111001110111000",
    "1111001110011111",
    "1111001111010010",
    "1111010001011001",
    "1111010100110001",
    "1111011001011000",
    "1111011111000010",
    "1111100101101001",
    "1111101101000000",
    "1111110101000101",
    "1111111101101110",
    "1111111001001010",
    "1111101111110110",
    "1111100110101000",
    "1111011101110011",
    "1111010101101100",
    "1111001110100001",
    "1111001000010110",
    "1111000011001101",
    "1110111110111011",
    "1110111011010110",
    "1110111000010001",
    "1110110101100100",
    "1110110011000101",
    "1110110000101100",
    "1110101110011100",
    "1110101100010111",
    "1110101010100000",
    "1110101000111100",
    "1110100111110010",
    "1110100111000100",
    "1110100110110111",
    "1110100111001000",
    "1110100111110100",
    "1110101000110111",
    "1110101010001100",
    "1110101011110010",
    "1110101101100110",
    "1110101111101011",
    "1110110010000010",
    "1110110100101110",
    "1110110111110100",
    "1110111011011000",
    "1110111111011010",
    "1111000011111100",
    "1111001000110111",
    "1111001110000000",
    "1111010011000110",
    "1111010111110010",
    "1111011011101000",
    "1111011110001111",
    "1111011111010111",
    "1111011110111101",
    "1111011101001010",
    "1111011010010011",
    "1111010110110010",
    "1111010011000101",
    "1111001111011110",
    "1111001100010011",
    "1111001001110000",
    "1111000111111111",
    "1111000111001001",
    "1111000111010101",
    "1111001000101101",
    "1111001011010110",
    "1111001111011100",
    "1111010101001001",
    "1111011100100110",
    "1111100101111011",
    "1111110001000000",
    "1111111101101001",
    "1111110100100111",
    "1111100110011111",
    "1111011000110100",
    "1111001100010111",
    "1111000001110001",
    "1110111001010101",
    "1110110011000000",
    "1110101110011001",
    "1110101010111000",
    "1110100111110010",
    "1110100100100100",
    "1110100000111000",
    "1110011100101110",
    "1110011000010000",
    "1110010011101110",
    "1110001111011001",
    "1110001011100001",
    "1110001000010011",
    "1110000101111001",
    "1110000100011101",
    "1110000100001011",
    "1110000101001101",
    "1110000111101000",
    "1110001011011110",
    "1110010000101110",
    "1110010111010101",
    "1110011111010010",
    "1110101000100010",
    "1110110010111110",
    "1110111110011011",
    "1111001010011001",
    "1111010110010011",
    "1111100001010000",
    "1111101010100000",
    "1111110001011001",
    "1111110101110000",
    "1111110111110100",
    "1111111000000101",
    "1111110111010000",
    "1111110101111110",
    "1111110100101010",
    "1111110011011111",
    "1111110010011100",
    "1111110001010101",
    "1111101111111111",
    "1111101110001011",
    "1111101011110000",
    "1111101000101101",
    "1111100101000110",
    "1111100001001100",
    "1111011101010100",
    "1111011001111010",
    "1111010111010110",
    "1111010101110110",
    "1111010101011111",
    "1111010110010010",
    "1111011000000100",
    "1111011010101111",
    "1111011110000101",
    "1111100001111110",
    "1111100110010011",
    "1111101010101110",
    "1111101111000001",
    "1111110010110100",
    "1111110101111001",
    "1111111000001011",
    "1111111001101100",
    "1111111010101001",
    "1111111011001101",
    "1111111011011110",
    "1111111011011001",
    "1111111010101101",
    "1111111001000011",
    "1111110110000010",
    "1111110001011011",
    "1111101011000111",
    "1111100011001111",
    "1111011010000110",
    "1111010000001000",
    "1111000101110110",
    "1110111011110011",
    "1110110010100111",
    "1110101010110101",
    "1110100100111100",
    "1110100001010000",
    "1110011111110000",
    "1110100000001111",
    "1110100010010000",
    "1110100101011101",
    "1110101001100101",
    "1110101110100001",
    "1110110100010111",
    "1110111011001001",
    "1111000010111001",
    "1111001011100001",
    "1111010100101100",
    "1111011101111111",
    "1111100110111000",
    "1111101110111011",
    "1111110101101011",
    "1111111010110101",
    "1111111110010001",
    "1111111111111001",
    "1111111111011110",
    "1111111111111001",
    "1111111110101101",
    "1111111101010011",
    "1111111011110110",
    "1111111010011000",
    "1111111000110010",
    "1111110110111011",
    "1111110100101001",
    "1111110001110110",
    "1111101110100101",
    "1111101010111010",
    "1111100110111110",
    "1111100010111101",
    "1111011111000010",
    "1111011011100011",
    "1111011000101111",
    "1111010110110001",
    "1111010101101100",
    "1111010101010101",
    "1111010101011010",
    "1111010101100100",
    "1111010101100010",
    "1111010101001110",
    "1111010100110111",
    "1111010100111001",
    "1111010101110110",
    "1111011000010001",
    "1111011100100110",
    "1111100010111011",
    "1111101011000001",
    "1111110100010111",
    "1111111110001100",
    "1111111000010010",
    "1111101111110101",
    "1111101000111110",
    "1111100011111100",
    "1111100000110110",
    "1111011111100110",
    "1111100000000010",
    "1111100010000110",
    "1111100101110010",
    "1111101011001100",
    "1111110010010110",
    "1111111011000110",
    "1111111011000000",
    "1111110000110010",
    "1111100111001000",
    "1111011110111000",
    "1111011000100111",
    "1111010100011100",
    "1111010010000101",
    "1111010001000010",
    "1111010000101011",
    "1111010000100110",
    "1111010000100100",
    "1111010000101100",
    "1111010001001010",
    "1111010010001111",
    "1111010100000001",
    "1111010110101000",
    "1111011001111100",
    "1111011101110101",
    "1111100010000110",
    "1111100110101010",
    "1111101011011100",
    "1111110000010110",
    "1111110101011011",
    "1111111010101000",
    "1111111111111101",
    "1111111010100100",
    "1111110101000100",
    "1111101111100111",
    "1111101010011000",
    "1111100101101100",
    "1111100001110110",
    "1111011111010001",
    "1111011110001010",
    "1111011110101001",
    "1111100000101001",
    "1111100011101111",
    "1111100111011111",
    "1111101011010100",
    "1111101110110000",
    "1111110001100000",
    "1111110011100001",
    "1111110100111101",
    "1111110110000011",
    "1111110111001000",
    "1111111000011011",
    "1111111010000011",
    "1111111011111110",
    "1111111110000001",
    "1111111111111001",
    "1111111110101011",
    "1111111110000001",
    "1111111110001010",
    "1111111111001001",
    "1111111111000110",
    "1111111100110011",
    "1111111010000011",
    "1111110110111110",
    "1111110011101001",
    "1111110000000100",
    "1111101100001100",
    "1111100111111110",
    "1111100011010011",
    "1111011110001101",
    "1111011000101000",
    "1111010010101001",
    "1111001100010001",
    "1111000101011011",
    "1110111110000111",
    "1110110110011010",
    "1110101110110001",
    "1110100111111001",
    "1110100010101001",
    "1110011111110011",
    "1110011111110000",
    "1110100010010000",
    "1110100110101010",
    "1110101011111000",
    "1110110000111101",
    "1110110101000001",
    "1110110111101100",
    "1110111000101111",
    "1110111000001011",
    "1110110110000000",
    "1110110010010000",
    "1110101101001010",
    "1110100110111011",
    "1110011111111011",
    "1110011000100111",
    "1110010001011001",
    "1110001010101010",
    "1110000100101010",
    "1101111111110000",
    "1101111100000111",
    "1101111010000001",
    "1101111001100011",
    "1101111010111000",
    "1101111110000101",
    "1110000011010000",
    "1110001010100010",
    "1110010011111110",
    "1110011111010111",
    "1110101100010001",
    "1110111001110100",
    "1111000111000100",
    "1111010011001010",
    "1111011101011001",
    "1111100101011111",
    "1111101011100101",
    "1111101111111110",
    "1111110011001100",
    "1111110101101110",
    "1111110111111111",
    "1111111010011010",
    "1111111101010000",
    "1111111111010000",
    "1111111011001001",
    "1111110110011100",
    "1111110001010101",
    "1111101100001010",
    "1111100111001110",
    "1111100010110110",
    "1111011111001010",
    "1111011100001110",
    "1111011001111010",
    "1111011000001001",
    "1111010110110001",
    "1111010101101110",
    "1111010101000101",
    "1111010100111110",
    "1111010101100100",
    "1111010111000001",
    "1111011001011101",
    "1111011100111010",
    "1111100001010010",
    "1111100110011100",
    "1111101100000101",
    "1111110001111010",
    "1111110111100000",
    "1111111100011111",
    "1111111111011100",
    "1111111100100011",
    "1111111010110110",
    "1111111010001111",
    "1111111010011101",
    "1111111011001111",
    "1111111100011000",
    "1111111101110010",
    "1111111111011011",
    "1111111110101001",
    "1111111100011110",
    "1111111001111101",
    "1111110111001101",
    "1111110100010000",
    "1111110001001110",
    "1111101110010100",
    "1111101011101010",
    "1111101001100010",
    "1111101000001010",
    "1111100111101111",
    "1111101000011101",
    "1111101010010111",
    "1111101101011101",
    "1111110001101000",
    "1111110110101101",
    "1111111100100001",
    "1111111101000010",
    "1111110110001001",
    "1111101110110000",
    "1111100110110011",
    "1111011110010100",
    "1111010101011011",
    "1111001100101000",
    "1111000100100111",
    "1110111110000101",
    "1110111001110000",
    "1110110111111100",
    "1110111000100010",
    "1110111011000110",
    "1110111110111101",
    "1111000011011101",
    "1111001000000011",
    "1111001100010100",
    "1111010000000101",
    "1111010011001011",
    "1111010101100101",
    "1111010111001000",
    "1111010111101010",
    "1111010110111111",
    "1111010101000000",
    "1111010001100110",
    "1111001100110011",
    "1111000110110111",
    "1111000000000111",
    "1110111000111110",
    "1110110010000010",
    "1110101011110101",
    "1110100110111001",
    "1110100011100001",
    "1110100001110110",
    "1110100001110000",
    "1110100011000000",
    "1110100101001101",
    "1110101000000001",
    "1110101011000010",
    "1110101110000000",
    "1110110000101110",
    "1110110011001000",
    "1110110101001101",
    "1110110111000110",
    "1110111001000001",
    "1110111011011000",
    "1110111110100100",
    "1111000011000011",
    "1111001001000110",
    "1111010000101011",
    "1111011001011110",
    "1111100010111011",
    "1111101100010100",
    "1111110101000001",
    "1111111100100111",
    "1111111101000111",
    "1111111000001110",
    "1111110100100011",
    "1111110001111001",
    "1111101111111111",
    "1111101110101010",
    "1111101101110101",
    "1111101101011010",
    "1111101101010110",
    "1111101101100100",
    "1111101101111011",
    "1111101110001100",
    "1111101110000100",
    "1111101101010011",
    "1111101011101010",
    "1111101001000011",
    "1111100101100010",
    "1111100001010100",
    "1111011100101000",
    "1111010111101101",
    "1111010010110011",
    "1111001110000000",
    "1111001001011110",
    "1111000101001110",
    "1111000001010010",
    "1110111101100001",
    "1110111001111001",
    "1110110110010011",
    "1110110010101110",
    "1110101111001010",
    "1110101011110010",
    "1110101000101100",
    "1110100110000000",
    "1110100011110100",
    "1110100010010100",
    "1110100001100100",
    "1110100001110011",
    "1110100011001000",
    "1110100101100101",
    "1110101001001001",
    "1110101101100011",
    "1110110010011010",
    "1110110111010101",
    "1110111011110101",
    "1110111111101011",
    "1111000010110001",
    "1111000101000101",
    "1111000110101101",
    "1111000111110100",
    "1111001000011101",
    "1111001000101010",
    "1111001000011101",
    "1111000111111100",
    "1111000111001011",
    "1111000110010010",
    "1111000101010111",
    "1111000100011000",
    "1111000011010101",
    "1111000010000010",
    "1111000000010100",
    "1110111110001001",
    "1110111011011110",
    "1110111000100000",
    "1110110101100000",
    "1110110010111011",
    "1110110001001000",
    "1110110000100001",
    "1110110001010010",
    "1110110011100010",
    "1110110111001011",
    "1110111011111101",
    "1111000001011010",
    "1111000110111111",
    "1111001100001010",
    "1111010000100001",
    "1111010011110011",
    "1111010101110110",
    "1111010110110100",
    "1111010110111001",
    "1111010110010010",
    "1111010101000110",
    "1111010011011000",
    "1111010001000101",
    "1111001110001001",
    "1111001010101010",
    "1111000110110110",
    "1111000010111110",
    "1110111111011111",
    "1110111100101101",
    "1110111010111000",
    "1110111010000111",
    "1110111010010100",
    "1110111011011011",
    "1110111101001111",
    "1110111111101110",
    "1111000010101110",
    "1111000110000110",
    "1111001001101101",
    "1111001101010001",
    "1111010000011110",
    "1111010010111110",
    "1111010100100000",
    "1111010100110110",
    "1111010011111100",
    "1111010001111001",
    "1111001110111101",
    "1111001011100000",
    "1111001000000001",
    "1111000101000001",
    "1111000011000001",
    "1111000010010111",
    "1111000011010000",
    "1111000101110110",
    "1111001010000110",
    "1111001111111101",
    "1111010111001110",
    "1111011111110000",
    "1111101001001111",
    "1111110011011000",
    "1111111101101111",
    "1111111000001110",
    "1111101111001100",
    "1111100111110010",
    "1111100010100111",
    "1111100000000111",
    "1111100000011001",
    "1111100011011010",
    "1111101000110111",
    "1111110000011011",
    "1111111001101101",
    "1111111011101000",
    "1111110000010001",
    "1111100100111001",
    "1111011010011011",
    "1111010001101110",
    "1111001011100000",
    "1111000111111111",
    "1111000111000100",
    "1111001000001110",
    "1111001010110100",
    "1111001110001101",
    "1111010010000101",
    "1111010110001000",
    "1111011010001110",
    "1111011110001100",
    "1111100001111011",
    "1111100101010010",
    "1111101000001111",
    "1111101010101110",
    "1111101100110010",
    "1111101110011010",
    "1111101111100100",
    "1111110000010100",
    "1111110000101100",
    "1111110000110001",
    "1111110000110000",
    "1111110000101111",
    "1111110000110101",
    "1111110001000001",
    "1111110001010101",
    "1111110001110001",
    "1111110010011000",
    "1111110011001100",
    "1111110100001111",
    "1111110101011110",
    "1111110110110100",
    "1111111000001110",
    "1111111001101000",
    "1111111011000101",
    "1111111100101100",
    "1111111110101001",
    "1111111110110110",
    "1111111011101000",
    "1111110111011011",
    "1111110010000111",
    "1111101011101101",
    "1111100100100000",
    "1111011101000111",
    "1111010110010011",
    "1111010000110011",
    "1111001101000010",
    "1111001011000010",
    "1111001010011000",
    "1111001010011110",
    "1111001010101010",
    "1111001010100000",
    "1111001001111001",
    "1111001000110101",
    "1111000111100000",
    "1111000101111100",
    "1111000100000110",
    "1111000001111110",
    "1110111111100011",
    "1110111101000010",
    "1110111010110000",
    "1110111001000100",
    "1110111000010110",
    "1110111000101010",
    "1110111001111101",
    "1110111100000001",
    "1110111110101000",
    "1111000001101110",
    "1111000101011011",
    "1111001001111111",
    "1111001111011111",
    "1111010101111100",
    "1111011101000010",
    "1111100100010011",
    "1111101011001111",
    "1111110001010101",
    "1111110110010011",
    "1111111010000111",
    "1111111100111010",
    "1111111110110100",
    "1111111111111010",
    "1111111111111000",
    "1111111111001011",
    "1111111101000100",
    "1111111001101111",
    "1111110101011000",
    "1111110000011000",
    "1111101011000101",
    "1111100101110010",
    "1111100000100011",
    "1111011011010001",
    "1111010101101111",
    "1111001111110001",
    "1111001001001011",
    "1111000001110000",
    "1110111001010110",
    "1110101111111000",
    "1110100101011101",
    "1110011010100101",
    "1110001111111011",
    "1110000110011111",
    "1101111111000111",
    "1101111010011000",
    "1101111000010011",
    "1101111000100000",
    "1101111010010110",
    "1101111101010010",
    "1110000000111110",
    "1110000101010111",
    "1110001010011110",
    "1110010000011010",
    "1110010111000100",
    "1110011110001100",
    "1110100101010011",
    "1110101100000010",
    "1110110010000011",
    "1110110111001000",
    "1110111011010001",
    "1110111110101000",
    "1111000001100001",
    "1111000100010011",
    "1111000111001110",
    "1111001010011011",
    "1111001101110010",
    "1111010001001100",
    "1111010100011010",
    "1111010111011011",
    "1111011010001111",
    "1111011100111111",
    "1111011111101011",
    "1111100010010000",
    "1111100100011111",
    "1111100110000100",
    "1111100110110010",
    "1111100110101010",
    "1111100110000011",
    "1111100101100000",
    "1111100101110001",
    "1111100111011001",
    "1111101010110001",
    "1111101111110101",
    "1111110110010000",
    "1111111101011101",
    "1111111011000010",
    "1111110011110001",
    "1111101100111111",
    "1111100110110100",
    "1111100001010000",
    "1111011100010011",
    "1111010111110111",
    "1111010100000000",
    "1111010000101011",
    "1111001101111101",
    "1111001011110101",
    "1111001010011000",
    "1111001001100000",
    "1111001001010101",
    "1111001001110010",
    "1111001010111010",
    "1111001100100110",
    "1111001110110011",
    "1111010001010101",
    "1111010100000101",
    "1111010110110010",
    "1111011001010101",
    "1111011011100001",
    "1111011101001111",
    "1111011110011100",
    "1111011111000100",
    "1111011111001000",
    "1111011110101101",
    "1111011101111000",
    "1111011100101110",
    "1111011011010110",
    "1111011001110000",
    "1111010111111111",
    "1111010110000100",
    "1111010011111110",
    "1111010001101100",
    "1111001111010010",
    "1111001100110000",
    "1111001010001111",
    "1111000111111100",
    "1111000110000110",
    "1111000101001001",
    "1111000101100111",
    "1111000111111100",
    "1111001100100000",
    "1111010011010010",
    "1111011011111101",
    "1111100101111011",
    "1111110000011001",
    "1111111010101010",
    "1111111011101110",
    "1111110011000011",
    "1111101011010110",
    "1111100100100111",
    "1111011110111010",
    "1111011010010001",
    "1111010110110111",
    "1111010100100101",
    "1111010011010000",
    "1111010010100001",
    "1111010001110100",
    "1111010000101011",
    "1111001110100110",
    "1111001011010001",
    "1111000110101101",
    "1111000001000010",
    "1110111010100101",
    "1110110011110011",
    "1110101101001100",
    "1110100111011000",
    "1110100010110001",
    "1110011111101110",
    "1110011110011011",
    "1110011110110011",
    "1110100000110000",
    "1110100011111001",
    "1110100111110111",
    "1110101100010100",
    "1110110000111011",
    "1110110101011101",
    "1110111001110101",
    "1110111110000100",
    "1111000010001000",
    "1111000110000110",
    "1111001001111101",
    "1111001101101001",
    "1111010001000000",
    "1111010011111000",
    "1111010110000110",
    "1111010111100111",
    "1111011000001110",
    "1111010111111001",
    "1111010110100000",
    "1111010100000011",
    "1111010000101001",
    "1111001100100011",
    "1111001000001011",
    "1111000011111110",
    "1111000000011100",
    "1110111101111101",
    "1110111100101101",
    "1110111100101010",
    "1110111101110010",
    "1111000000000000",
    "1111000011010010",
    "1111000111110001",
    "1111001101101001",
    "1111010101000110",
    "1111011110001010",
    "1111101000101110",
    "1111110100100011",
    "1111111110101011",
    "1111110001100010",
    "1111100100100000",
    "1111011000001110",
    "1111001101001111",
    "1111000100000000",
    "1110111100101000",
    "1110110110111110",
    "1110110010100111",
    "1110101110111111",
    "1110101011100000",
    "1110100111110001",
    "1110100011100100",
    "1110011110111000",
    "1110011001110101",
    "1110010100100101",
    "1110001111010111",
    "1110001010011011",
    "1110000110001101",
    "1110000011000110",
    "1110000001100100",
    "1110000001111101",
    "1110000100011000",
    "1110001000111010",
    "1110001111011110",
    "1110010111111001",
    "1110100001111001",
    "1110101101010001",
    "1110111001100111",
    "1111000110100000",
    "1111010011010101",
    "1111011111010010",
    "1111101001011111",
    "1111110001010100",
    "1111110110010111",
    "1111111000110000",
    "1111111001000000",
    "1111110111110110",
    "1111110110001000",
    "1111110100011001",
    "1111110010111110",
    "1111110001111001",
    "1111110001000011",
    "1111110000011010",
    "1111101111111100",
    "1111101111101110",
    "1111101111110010",
    "1111110000000111",
    "1111110000100111",
    "1111110001001011",
    "1111110001101011",
    "1111110010001001",
    "1111110010100110",
    "1111110011001000",
    "1111110011101101",
    "1111110100010001",
    "1111110100110001",
    "1111110101001010",
    "1111110101100010",
    "1111110101111100",
    "1111110110011101",
    "1111110111000011",
    "1111110111100101",
    "1111110111111110",
    "1111111000001001",
    "1111111000001100",
    "1111111000010010",
    "1111111000100001",
    "1111111000110101",
    "1111111000111011",
    "1111111000010100",
    "1111110110011100",
    "1111110010110110",
    "1111101101010010",
    "1111100101110001",
    "1111011100100101",
    "1111010010001011",
    "1111000111001110",
    "1110111100011001",
    "1110110010010111",
    "1110101001101111",
    "1110100011000001",
    "1110011110011100",
    "1110011100000001",
    "1110011011100000",
    "1110011100100101",
    "1110011110111011",
    "1110100010010010",
    "1110100110100000",
    "1110101011100000",
    "1110110001010100",
    "1110111000000001",
    "1110111111101011",
    "1111001000010000",
    "1111010001100111",
    "1111011011011011",
    "1111100101000101",
    "1111101101110110",
    "1111110100111011",
    "1111111001110011",
    "1111111100010111",
    "1111111100111011",
    "1111111100001101",
    "1111111011000000",
    "1111111010000000",
    "1111111001100010",
    "1111111001100011",
    "1111111001101010",
    "1111111001011000",
    "1111111000001110",
    "1111110101110110",
    "1111110010000110",
    "1111101100111011",
    "1111100110011001",
    "1111011110101001",
    "1111010110000001",
    "1111001101000010",
    "1111000100011100",
    "1110111101000010",
    "1110110111101000",
    "1110110100101110",
    "1110110100011010",
    "1110110110010110",
    "1110111001110111",
    "1110111110001101",
    "1111000010110011",
    "1111000111010110",
    "1111001011111101",
    "1111010001000000",
    "1111010110111100",
    "1111011110000010",
    "1111100110001101",
    "1111101111000101",
    "1111111000000111",
    "1111111111001100",
    "1111110111010111",
    "1111110000100101",
    "1111101011000110",
    "1111100110111111",
    "1111100100011101",
    "1111100011101010",
    "1111100100110100",
    "1111101000000101",
    "1111101101100011",
    "1111110101001111",
    "1111111110110100",
    "1111110110010001",
    "1111101011000010",
    "1111100000100110",
    "1111010111111001",
    "1111010001100001",
    "1111001101100011",
    "1111001011100001",
    "1111001010101010",
    "1111001010001011",
    "1111001001100111",
    "1111001000110100",
    "1111001000001000",
    "1111000111110111",
    "1111001000100010",
    "1111001010010011",
    "1111001101001100",
    "1111010001000011",
    "1111010101100111",
    "1111011010101101",
    "1111100000001000",
    "1111100101110010",
    "1111101011100110",
    "1111110001011100",
    "1111110111001100",
    "1111111100101111",
    "1111111101111101",
    "1111111001001000",
    "1111110100110011",
    "1111110001000110",
    "1111101110000110",
    "1111101011110001",
    "1111101010000000",
    "1111101000101000",
    "1111100111011100",
    "1111100110011001",
    "1111100101100000",
    "1111100100111110",
    "1111100101000001",
    "1111100101111001",
    "1111100111101011",
    "1111101010010101",
    "1111101101101010",
    "1111110001010110",
    "1111110101000111",
    "1111111000101000",
    "1111111011110000",
    "1111111110010000",
    "1111111111110110",
    "1111111110101001",
    "1111111110000100",
    "1111111101111101",
    "1111111110001111",
    "1111111110110101",
    "1111111111110000",
    "1111111110111010",
    "1111111101000111",
    "1111111010101110",
    "1111110111101111",
    "1111110100001100",
    "1111110000001011",
    "1111101011110111",
    "1111100111010111",
    "1111100010110100",
    "1111011110010001",
    "1111011001101101",
    "1111010100110110",
    "1111001111011001",
    "1111001000111001",
    "1111000001001101",
    "1110111000100011",
    "1110101111101001",
    "1110100111011011",
    "1110100000111001",
    "1110011100110011",
    "1110011011011110",
    "1110011100101101",
    "1110011111111101",
    "1110100100100111",
    "1110101010000010",
    "1110101111101001",
    "1110110100110011",
    "1110111000110100",
    "1110111010111101",
    "1110111010100110",
    "1110110111010110",
    "1110110001001101",
    "1110101000100111",
    "1110011110011001",
    "1110010011100100",
    "1110001001000110",
    "1101111111110101",
    "1101111000010001",
    "1101110010101111",
    "1101101111010100",
    "1101101101111111",
    "1101101110101101",
    "1101110001011111",
    "1101110110011010",
    "1101111101011100",
    "1110000110011101",
    "1110010001000011",
    "1110011100100101",
    "1110101000011000",
    "1110110011101110",
    "1110111110001001",
    "1111000111010110",
    "1111001111011001",
    "1111010110010010",
    "1111011100000111",
    "1111100000111011",
    "1111100100101111",
    "1111100111101101",
    "1111101010000110",
    "1111101100010100",
    "1111101110111001",
    "1111110010010010",
    "1111110110110111",
    "1111111100101001",
    "1111111100100011",
    "1111110101010010",
    "1111101110001000",
    "1111100111101001",
    "1111100010010100",
    "1111011110011001",
    "1111011011111100",
    "1111011010111010",
    "1111011011000110",
    "1111011100010100",
    "1111011110010111",
    "1111100001000111",
    "1111100100011010",
    "1111101000001110",
    "1111101100011001",
    "1111110000110110",
    "1111110101011010",
    "1111111001111000",
    "1111111110000010",
    "1111111110010100",
    "1111111011011100",
    "1111111001011001",
    "1111111000001111",
    "1111110111111001",
    "1111111000001100",
    "1111111000111011",
    "1111111001111001",
    "1111111011000000",
    "1111111100010001",
    "1111111101110110",
    "1111111111111010",
    "1111111101010110",
    "1111111001111100",
    "1111110101111001",
    "1111110001011101",
    "1111101100111100",
    "1111101000101111",
    "1111100101010000",
    "1111100010101111",
    "1111100001011110",
    "1111100001011111",
    "1111100010110011",
    "1111100101010101",
    "1111101000111110",
    "1111101101100110",
    "1111110011000111",
    "1111111001010101",
    "1111111111111001",
    "1111111000110011",
    "1111110001101001",
    "1111101010100111",
    "1111100011111001",
    "1111011101100110",
    "1111010111110100",
    "1111010010110001",
    "1111001110101101",
    "1111001011111000",
    "1111001010011110",
    "1111001010011110",
    "1111001011101000",
    "1111001101100110",
    "1111001111111010",
    "1111010010001010",
    "1111010100000011",
    "1111010101010111",
    "1111010110000000",
    "1111010110000000",
    "1111010101011101",
    "1111010100100010",
    "1111010011011100",
    "1111010010010111",
    "1111010001010101",
    "1111010000001111",
    "1111001110110000",
    "1111001100100001",
    "1111001001010110",
    "1111000101001101",
    "1111000000010001",
    "1110111010111100",
    "1110110101110100",
    "1110110001010100",
    "1110101101110101",
    "1110101011100101",
    "1110101010100110",
    "1110101010110111",
    "1110101100001010",
    "1110101110010110",
    "1110110001001000",
    "1110110100010011",
    "1110110111101100",
    "1110111011001010",
    "1110111110101101",
    "1111000010001111",
    "1111000101110001",
    "1111001001010110",
    "1111001101000000",
    "1111010000111000",
    "1111010101000101",
    "1111011001101111",
    "1111011110111101",
    "1111100100101110",
    "1111101010110111",
    "1111110001001100",
    "1111110111011011",
    "1111111101010111",
    "1111111101000101",
    "1111111000000010",
    "1111110011011101",
    "1111101111011000",
    "1111101011110101",
    "1111101000111100",
    "1111100110110010",
    "1111100101010111",
    "1111100100100101",
    "1111100100010010",
    "1111100100010000",
    "1111100100010010",
    "1111100100001011",
    "1111100011101010",
    "1111100010100111",
    "1111100000111011",
    "1111011110100001",
    "1111011011011011",
    "1111010111110010",
    "1111010011101110",
    "1111001111010110",
    "1111001010101101",
    "1111000101110111",
    "1111000000111001",
    "1110111011111000",
    "1110110110111110",
    "1110110010011001",
    "1110101110010110",
    "1110101011000001",
    "1110101000100101",
    "1110100111010000",
    "1110100111001000",
    "1110101000010001",
    "1110101010101101",
    "1110101110001001",
    "1110110010001101",
    "1110110110011000",
    "1110111010000110",
    "1110111100111010",
    "1110111110100100",
    "1110111111000111",
    "1110111110111000",
    "1110111110010010",
    "1110111101111010",
    "1110111110000111",
    "1110111111000111",
    "1111000000110001",
    "1111000010110011",
    "1111000100110011",
    "1111000110100000",
    "1111000111110100",
    "1111001000101111",
    "1111001001010011",
    "1111001001011011",
    "1111001000111100",
    "1111000111100011",
    "1111000101000001",
    "1111000001010010",
    "1110111100100101",
    "1110110111011010",
    "1110110010010111",
    "1110101110000101",
    "1110101010111100",
    "1110101001001100",
    "1110101001000001",
    "1110101010100000",
    "1110101101101110",
    "1110110010101110",
    "1110111001010101",
    "1111000001001100",
    "1111001001101010",
    "1111010001111110",
    "1111011001010101",
    "1111011111001000",
    "1111100011000101",
    "1111100101001001",
    "1111100101011101",
    "1111100100001110",
    "1111100001100111",
    "1111011101101101",
    "1111011000100000",
    "1111010010001011",
    "1111001011000001",
    "1111000011101001",
    "1110111100110101",
    "1110110111011101",
    "1110110100010000",
    "1110110011101001",
    "1110110101101001",
    "1110111001111001",
    "1110111111110011",
    "1111000110100101",
    "1111001101100000",
    "1111010011110110",
    "1111011001000110",
    "1111011100110010",
    "1111011110100100",
    "1111011110010100",
    "1111011100000010",
    "1111010111111111",
    "1111010010100100",
    "1111001100010100",
    "1111000101110111",
    "1110111111110110",
    "1110111010110010",
    "1110110111001000",
    "1110110101001101",
    "1110110101010101",
    "1110110111110010",
    "1110111100100110",
    "1111000011101111",
    "1111001100110011",
    "1111010111010001",
    "1111100010011101",
    "1111101101100111",
    "1111111000001011",
    "1111111110010010",
    "1111110110001010",
    "1111101111100111",
    "1111101010110010",
    "1111100111110010",
    "1111100110100111",
    "1111100111001011",
    "1111101001001111",
    "1111101100100100",
    "1111110000111000",
    "1111110101111101",
    "1111111011100110",
    "1111111110010000",
    "1111110111111000",
    "1111110001011111",
    "1111101011011100",
    "1111100110001001",
    "1111100010000101",
    "1111011111100110",
    "1111011110111000",
    "1111011111111010",
    "1111100010011001",
    "1111100101110100",
    "1111101001100110",
    "1111101101000111",
    "1111101111111001",
    "1111110001110010",
    "1111110010110000",
    "1111110010111110",
    "1111110010100100",
    "1111110001101011",
    "1111110000010101",
    "1111101110101000",
    "1111101100101010",
    "1111101010101100",
    "1111101000111111",
    "1111100111101100",
    "1111100110111000",
    "1111100110011011",
    "1111100110001001",
    "1111100101111001",
    "1111100101101001",
    "1111100101011010",
    "1111100101010111",
    "1111100101101001",
    "1111100110010011",
    "1111100111011000",
    "1111101000110101",
    "1111101010100110",
    "1111101100101010",
    "1111101111000011",
    "1111110001110001",
    "1111110100111001",
    "1111111000011111",
    "1111111100101011",
    "1111111110011101",
    "1111111000111010",
    "1111110010110000",
    "1111101100001010",
    "1111100101011011",
    "1111011110111101",
    "1111011000111111",
    "1111010011101100",
    "1111001111000100",
    "1111001010111100",
    "1111000111001001",
    "1111000011100110",
    "1111000000010010",
    "1110111101010110",
    "1110111010111101",
    "1110111001010011",
    "1110111000100010",
    "1110111000101111",
    "1110111010000001",
    "1110111100010100",
    "1110111111100100",
    "1111000011011101",
    "1111000111100010",
    "1111001011010110",
    "1111001110011111",
    "1111010000110001",
    "1111010010010000",
    "1111010011010111",
    "1111010100100010",
    "1111010110011010",
    "1111011001011001",
    "1111011101110010",
    "1111100011011100",
    "1111101010000111",
    "1111110001010101",
    "1111111000101011",
    "1111111111101100",
    "1111111001111010",
    "1111110100011101",
    "1111110000000111",
    "1111101101000100",
    "1111101011011110",
    "1111101011011101",
    "1111101100111111",
    "1111101111111110",
    "1111110100001100",
    "1111111001011010",
    "1111111111011100",
    "1111111001110110",
    "1111110010101011",
    "1111101011000111",
    "1111100011010011",
    "1111011011011011",
    "1111010011101110",
    "1111001100010001",
    "1111000101001011",
    "1110111110011100",
    "1110111000000001",
    "1110110001110001",
    "1110101011101111",
    "1110100101111001",
    "1110100000011001",
    "1110011011011000",
    "1110010110111111",
    "1110010011011100",
    "1110010000110001",
    "1110001111000111",
    "1110001110010110",
    "1110001110010111",
    "1110001111000010",
    "1110010000010010",
    "1110010010000011",
    "1110010100011100",
    "1110010111011111",
    "1110011011010100",
    "1110011111111010",
    "1110100101001000",
    "1110101010110111",
    "1110110000111000",
    "1110110110111011",
    "1110111100101011",
    "1111000001111000",
    "1111000110001011",
    "1111001001010110",
    "1111001011010100",
    "1111001100001010",
    "1111001100001010",
    "1111001011101010",
    "1111001011000001",
    "1111001010101000",
    "1111001010101111",
    "1111001011100011",
    "1111001101001111",
    "1111001111110110",
    "1111010011010101",
    "1111010111100000",
    "1111011100001001",
    "1111100001000010",
    "1111100110000000",
    "1111101010111101",
    "1111101111111100",
    "1111110101000000",
    "1111111010001011",
    "1111111111010110",
    "1111111011101010",
    "1111110111001000",
    "1111110011001011",
    "1111101111110000",
    "1111101100101011",
    "1111101001101010",
    "1111100110011100",
    "1111100010110110",
    "1111011110111010",
    "1111011010110100",
    "1111010110110110",
    "1111010011010011",
    "1111010000011110",
    "1111001110100001",
    "1111001101101000",
    "1111001101110101",
    "1111001111001111",
    "1111010001110001",
    "1111010101010101",
    "1111011001101010",
    "1111011110011001",
    "1111100011000110",
    "1111100111010111",
    "1111101010101111",
    "1111101100111011",
    "1111101101101101",
    "1111101101000010",
    "1111101011000011",
    "1111101000000000",
    "1111100100010010",
    "1111100000010010",
    "1111011100011100",
    "1111011000111111",
    "1111010110001001",
    "1111010011111011",
    "1111010010001101",
    "1111010000111101",
    "1111010000000010",
    "1111001111011111",
    "1111001111011001",
    "1111001111111010",
    "1111010001001100",
    "1111010011011101",
    "1111010110110100",
    "1111011011000111",
    "1111100000001101",
    "1111100101110001",
    "1111101011011011",
    "1111110000111000",
    "1111110110000001",
    "1111111010110010",
    "1111111111001101",
    "1111111100101000",
    "1111111000110010",
    "1111110101010101",
    "1111110010010111",
    "1111101111111100",
    "1111101110000011",
    "1111101100011111",
    "1111101010110110",
    "1111101000100110",
    "1111100101001110",
    "1111100000010111",
    "1111011001110111",
    "1111010001111011",
    "1111001000111111",
    "1110111111101110",
    "1110110110110100",
    "1110101110111011",
    "1110101000011101",
    "1110100011101010",
    "1110100000101001",
    "1110011111010110",
    "1110011111100100",
    "1110100001001000",
    "1110100011101001",
    "1110100110101100",
    "1110101001110100",
    "1110101100100101",
    "1110101110110001",
    "1110110000010101",
    "1110110001100110",
    "1110110010111110",
    "1110110100111110",
    "1110110111101101",
    "1110111011000111",
    "1110111110101011",
    "1111000001110001",
    "1111000011110110",
    "1111000100100000",
    "1111000011101110",
    "1111000001101100",
    "1110111110110001",
    "1110111011011110",
    "1110111000001001",
    "1110110101001011",
    "1110110010111000",
    "1110110001011110",
    "1110110001000101",
    "1110110001110001",
    "1110110011011010",
    "1110110101111011",
    "1110111001000111",
    "1110111100111010",
    "1111000001010010",
    "1111000110010011",
    "1111001100000010",
    "1111010010100100",
    "1111011001110111",
    "1111100001110100",
    "1111101010010001",
    "1111110011000001",
    "1111111011111100",
    "1111111011000010",
    "1111110010000100",
    "1111101001000110",
    "1111100000000111",
    "1111010111001001",
    "1111001110001101",
    "1111000101010111",
    "1110111100101010",
    "1110110100001011",
    "1110101100000010",
    "1110100100010111",
    "1110011101010110",
    "1110010111001101",
    "1110010010001101",
    "1110001110100110",
    "1110001100100000",
    "1110001011111100",
    "1110001100110011",
    "1110001111000000",
    "1110010010011010",
    "1110010110111011",
    "1110011100011001",
    "1110100010101011",
    "1110101001100000",
    "1110110000101100",
    "1110111000000100",
    "1110111111011110",
    "1111000110110100",
    "1111001110000000",
    "1111010100110110",
    "1111011010111111",
    "1111100000000010",
    "1111100011101110",
    "1111100101111110",
    "1111100110111010",
    "1111100110110111",
    "1111100110010000",
    "1111100101011101",
    "1111100100110001",
    "1111100100010010",
    "1111100100000011",
    "1111100100000110",
    "1111100100011000",
    "1111100100110110",
    "1111100101011000",
    "1111100101111011",
    "1111100110010101",
    "1111100110100011",
    "1111100110100001",
    "1111100110010011",
    "1111100101111110",
    "1111100101110001",
    "1111100101111011",
    "1111100110101111",
    "1111101000011101",
    "1111101011001111",
    "1111101110111100",
    "1111110011010001",
    "1111110111100100",
    "1111111011001011",
    "1111111101011110",
    "1111111110000110",
    "1111111100111110",
    "1111111010011010",
    "1111110110110111",
    "1111110010110000",
    "1111101110011101",
    "1111101010000111",
    "1111100101101100",
    "1111100001000101",
    "1111011100000111",
    "1111010110110001",
    "1111010000111101",
    "1111001010110000",
    "1111000100001101",
    "1110111101010111",
    "1110110110010101",
    "1110101111010010",
    "1110101000011110",
    "1110100010010100",
    "1110011101000111",
    "1110011001001110",
    "1110010110110110",
    "1110010110000011",
    "1110010110101101",
    "1110011000110000",
    "1110011011111101",
    "1110100000001111",
    "1110100101100111",
    "1110101100001010",
    "1110110100000000",
    "1110111101000111",
    "1111000111010001",
    "1111010010000010",
    "1111011100101010",
    "1111100110011100",
    "1111101110101110",
    "1111110101000101",
    "1111111001011101",
    "1111111100000100",
    "1111111101010001",
    "1111111101011111",
    "1111111100111111",
    "1111111011111100",
    "1111111010010111",
    "1111111000001000",
    "1111110101001110",
    "1111110001100110",
    "1111101101010111",
    "1111101000101010",
    "1111100011101001",
    "1111011110010111",
    "1111011000111010",
    "1111010011010011",
    "1111001101100100",
    "1111000111111010",
    "1111000010101011",
    "1110111110001001",
    "1110111010100110",
    "1110111000001110",
    "1110110110111111",
    "1110110110110010",
    "1110110111100000",
    "1110111001000111",
    "1110111011101011",
    "1110111111011001",
    "1111000100011111",
    "1111001011001100",
    "1111010011101010",
    "1111011101111011",
    "1111101001101101",
    "1111110110011101",
    "1111111100101010",
    "1111110000110000",
    "1111100110101111",
    "1111011111010010",
    "1111011010110000",
    "1111011001000100",
    "1111011001110111",
    "1111011100110010",
    "1111100001100001",
    "1111100111111111",
    "1111110000001001",
    "1111111001111000",
    "1111111011001010",
    "1111101111101110",
    "1111100100101110",
    "1111011011000110",
    "1111010011100100",
    "1111001110100011",
    "1111001011110111",
    "1111001011000110",
    "1111001011100110",
    "1111001100110010",
    "1111001110001010",
    "1111001111100001",
    "1111010000110101",
    "1111010010001010",
    "1111010011101010",
    "1111010101011101",
    "1111010111101010",
    "1111011010010110",
    "1111011101100001",
    "1111100001010010",
    "1111100101101001",
    "1111101010100010",
    "1111101111110011",
    "1111110101001111",
    "1111111010100001",
    "1111111111010110",
    "1111111100011110",
    "1111111001001000",
    "1111110110100111",
    "1111110100110010",
    "1111110011011111",
    "1111110010011110",
    "1111110001100000",
    "1111110000011001",
    "1111101111000001",
    "1111101101010100",
    "1111101011010100",
    "1111101001000110",
    "1111100110110101",
    "1111100100110001",
    "1111100011001101",
    "1111100010011010",
    "1111100010100110",
    "1111100011111000",
    "1111100110010000",
    "1111101001101100",
    "1111101110000000",
    "1111110010110111",
    "1111110111111000",
    "1111111100100001",
    "1111111111101011",
    "1111111101001110",
    "1111111100010010",
    "1111111100110111",
    "1111111110110000",
    "1111111110010001",
    "1111111010100011",
    "1111110110001100",
    "1111110001010011",
    "1111101011110110",
    "1111100101111011",
    "1111011111100110",
    "1111011001000010",
    "1111010010011100",
    "1111001011111101",
    "1111000101110110",
    "1111000000010001",
    "1110111011011110",
    "1110110111101111",
    "1110110101010000",
    "1110110100000110",
    "1110110100010000",
    "1110110101100010",
    "1110110111101000",
    "1110111010001100",
    "1110111100110000",
    "1110111110111011",
    "1111000000010111",
    "1111000000110000",
    "1110111111111010",
    "1110111101110011",
    "1110111010011101",
    "1110110101111110",
    "1110110000100011",
    "1110101010011000",
    "1110100011101111",
    "1110011100111010",
    "1110010110001001",
    "1110001111101100",
    "1110001001110100",
    "1110000100100101",
    "1110000000001100",
    "1101111100100110",
    "1101111001111010",
    "1101111000001011",
    "1101110111011000",
    "1101110111100011",
    "1101111000101010",
    "1101111010101010",
    "1101111101100001",
    "1110000001001100",
    "1110000101101010",
    "1110001011000010",
    "1110010001010100",
    "1110011000100011",
    "1110100000110011",
    "1110101001111101",
    "1110110011110011",
    "1110111101111101",
    "1111001000001000",
    "1111010001110110",
    "1111011010111100",
    "1111100011010000",
    "1111101010110110",
    "1111110001111000",
    "1111111000100000",
    "1111111110110110",
    "1111111011000001",
    "1111110101010010",
    "1111110000000000",
    "1111101011001110",
    "1111100110111011",
    "1111100011000001",
    "1111011111011010",
    "1111011100000001",
    "1111011000111001",
    "1111010110010010",
    "1111010100011111",
    "1111010011110100",
    "1111010100100100",
    "1111010110101111",
    "1111011010010011",
    "1111011111000010",
    "1111100100101010",
    "1111101010110110",
    "1111110001001110",
    "1111110111010111",
    "1111111100110100",
    "1111111110110101",
    "1111111100000100",
    "1111111011000010",
    "1111111011101111",
    "1111111101111000",
    "1111111110111111",
    "1111111011011101",
    "1111110111111110",
    "1111110100110111",
    "1111110010010010",
    "1111110000001001",
    "1111101110010001",
    "1111101100011010",
    "1111101010011011",
    "1111101000010000",
    "1111100110000000",
    "1111100011111000",
    "1111100010001010",
    "1111100001000111",
    "1111100000111101",
    "1111100001110000",
    "1111100011100010",
    "1111100110010011",
    "1111101001111101",
    "1111101110011011",
    "1111110011100000",
    "1111111001000001",
    "1111111110101100",
    "1111111011101101",
    "1111110110011110",
    "1111110001101100",
    "1111101101010111",
    "1111101001011011",
    "1111100101110100",
    "1111100010100110",
    "1111011111101110",
    "1111011101010100",
    "1111011011011101",
    "1111011010001100",
    "1111011001100111",
    "1111011001110010",
    "1111011010110000",
    "1111011100100001",
    "1111011110110101",
    "1111100001011001",
    "1111100011101100",
    "1111100101001110",
    "1111100101101001",
    "1111100100101100",
    "1111100010010101",
    "1111011110101011",
    "1111011010000001",
    "1111010100101001",
    "1111001110111010",
    "1111001001000100",
    "1111000011010111",
    "1110111101111101",
    "1110111000111110",
    "1110110100011111",
    "1110110000100111",
    "1110101101100100",
    "1110101011011101",
    "1110101010011011",
    "1110101010100011",
    "1110101011110000",
    "1110101101110111",
    "1110110000100111",
    "1110110011101111",
    "1110110110111100",
    "1110111001111111",
    "1110111100101101",
    "1110111111000010",
    "1111000000111011",
    "1111000010011100",
    "1111000011101110",
    "1111000101000000",
    "1111000110100100",
    "1111001000101101",
    "1111001011100101",
    "1111001111010001",
    "1111010011100111",
    "1111011000011101",
    "1111011101100001",
    "1111100010101011",
    "1111100111110001",
    "1111101100110100",
    "1111110001110100",
    "1111110110110000",
    "1111111011011110",
    "1111111111110111",
    "1111111100001110",
    "1111111001000000",
    "1111110110011110",
    "1111110100100100",
    "1111110011000111",
    "1111110001110100",
    "1111110000011100",
    "1111101110110000",
    "1111101100101001",
    "1111101010000101",
    "1111100111001001",
    "1111100011111001",
    "1111100000011001",
    "1111011100101010",
    "1111011000101010",
    "1111010100011101",
    "1111010000001100",
    "1111001011111101",
    "1111000111111100",
    "1111000100010010",
    "1111000000111011",
    "1110111101110011",
    "1110111010110000",
    "1110110111101000",
    "1110110100011101",
    "1110110001010010",
    "1110101110010010",
    "1110101011101011",
    "1110101001101111",
    "1110101000101000",
    "1110101000011101",
    "1110101001010000",
    "1110101011000010",
    "1110101101110010",
    "1110110001010101",
    "1110110101101001",
    "1110111010011011",
    "1110111111011100",
    "1111000100010111",
    "1111001000110101",
    "1111001100101000",
    "1111001111100100",
    "1111010001100110",
    "1111010010110100",
    "1111010011010010",
    "1111010011000001",
    "1111010010000101",
    "1111010000011100",
    "1111001110000101",
    "1111001011001100",
    "1111001000000011",
    "1111000101000011",
    "1111000010100110",
    "1111000000111101",
    "1111000000010101",
    "1111000000100111",
    "1111000001100111",
    "1111000011001010",
    "1111000100111110",
    "1111000111000001",
    "1111001001001110",
    "1111001011101010",
    "1111001110010010",
    "1111010001000111",
    "1111010011111011",
    "1111010110100100",
    "1111011000101111",
    "1111011010010001",
    "1111011011000010",
    "1111011011000100",
    "1111011010011001",
    "1111011001001001",
    "1111010111011000",
    "1111010101000110",
    "1111010010010100",
    "1111001110111011",
    "1111001011000100",
    "1111000110111100",
    "1111000010111101",
    "1110111111100011",
    "1110111101001110",
    "1110111100010001",
    "1110111100110101",
    "1110111110110001",
    "1111000001110001",
    "1111000101011011",
    "1111001001001110",
    "1111001100101110",
    "1111001111100001",
    "1111010001010111",
    "1111010010000101",
    "1111010001101100",
    "1111010000010111",
    "1111001110010100",
    "1111001011110101",
    "1111001001010000",
    "1111000110110010",
    "1111000100100111",
    "1111000010111000",
    "1111000001101001",
    "1111000001000011",
    "1111000001010010",
    "1111000010100001",
    "1111000100110110",
    "1111001000011000",
    "1111001101000100",
    "1111010010110100",
    "1111011001100000",
    "1111100000110110",
    "1111101000100010",
    "1111110000000010",
    "1111110110111001",
    "1111111100100100",
    "1111111111001111",
    "1111111100110010",
    "1111111100000010",
    "1111111100111000",
    "1111111111001011",
    "1111111101001000",
    "1111111000010000",
    "1111110010010010",
    "1111101011100101",
    "1111100100100100",
    "1111011101111000",
    "1111011000001100",
    "1111010100001010",
    "1111010010001000",
    "1111010010010100",
    "1111010100100100",
    "1111011000101000",
    "1111011110000010",
    "1111100100001010",
    "1111101010010111",
    "1111101111111110",
    "1111110100011011",
    "1111110111010010",
    "1111111000010100",
    "1111110111100011",
    "1111110101001011",
    "1111110001101001",
    "1111101101011011",
    "1111101001000011",
    "1111100100111100",
    "1111100001010111",
    "1111011110011110",
    "1111011100001111",
    "1111011010101101",
    "1111011001101111",
    "1111011001010101",
    "1111011001011001",
    "1111011001110111",
    "1111011010100101",
    "1111011011010110",
    "1111011100000100",
    "1111011100100110",
    "1111011100111010",
    "1111011101000101",
    "1111011101001110",
    "1111011101011100",
    "1111011101111000",
    "1111011110101101",
    "1111100000000000",
    "1111100001111101",
    "1111100100101010",
    "1111101000010010",
    "1111101100111011",
    "1111110010101001",
    "1111111001011111",
    "1111111110100001",
    "1111110101100011",
    "1111101011111010",
    "1111100010001101",
    "1111011001001100",
    "1111010001101100",
    "1111001100010100",
    "1111001001001110",
    "1111001000001110",
    "1111001000101000",
    "1111001001101010",
    "1111001010100010",
    "1111001010101101",
    "1111001010000010",
    "1111001000100010",
    "1111000110100000",
    "1111000100010000",
    "1111000010000101",
    "1111000000001101",
    "1110111110101110",
    "1110111101110010",
    "1110111101010110",
    "1110111101100000",
    "1110111110001111",
    "1110111111101110",
    "1111000010010000",
    "1111000110000110",
    "1111001011100101",
    "1111010010111000",
    "1111011011110010",
    "1111100101110110",
    "1111110000010000",
    "1111111010001100",
    "1111111100111110",
    "1111110101110010",
    "1111110000011010",
    "1111101100110110",
    "1111101011000001",
    "1111101010110011",
    "1111101100000011",
    "1111101110101000",
    "1111110010010011",
    "1111110110110010",
    "1111111011101111",
    "1111111111000110",
    "1111111001111111",
    "1111110100111101",
    "1111101111111110",
    "1111101010110111",
    "1111100101100010",
    "1111011111110101",
    "1111011001101010",
    "1111010011000000",
    "1111001011110101",
    "1111000100000110",
    "1110111011111101",
    "1110110011011101",
    "1110101010111101",
    "1110100010110011",
    "1110011011011101",
    "1110010101011000",
    "1110010000111001",
    "1110001110001010",
    "1110001101000010",
    "1110001101001110",
    "1110001110001101",
    "1110001111101001",
    "1110010001001111",
    "1110010010110011",
    "1110010100010111",
    "1110010110000000",
    "1110010111110010",
    "1110011001110000",
    "1110011011111101",
    "1110011110011011",
    "1110100001010100",
    "1110100100101110",
    "1110101000110101",
    "1110101101101101",
    "1110110011001011",
    "1110111001000010",
    "1110111110111010",
    "1111000100010111",
    "1111001001000010",
    "1111001100101110",
    "1111001111010111",
    "1111010001000010",
    "1111010001110110",
    "1111010010000101",
    "1111010001111001",
    "1111010001100010",
    "1111010001001000",
    "1111010000110101",
    "1111010000110000",
    "1111010001000011",
    "1111010010000000",
    "1111010011101110",
    "1111010110011010",
    "1111011001111101",
    "1111011110001111",
    "1111100010111000",
    "1111100111100010",
    "1111101011111001",
    "1111101111110101",
    "1111110011011011",
    "1111110110110111",
    "1111111010011011",
    "1111111110011001",
    "1111111101000101",
    "1111111000001000",
    "1111110010111011",
    "1111101101110011",
    "1111101001001000",
    "1111100101010000",
    "1111100010011010",
    "1111100000101001",
    "1111011111111011",
    "1111100000000000",
    "1111100000100111",
    "1111100001100010",
    "1111100010100100",
    "1111100011100111",
    "1111100100101001",
    "1111100101100101",
    "1111100110011001",
    "1111100110111001",
    "1111100110111010",
    "1111100110010010",
    "1111100100111001",
    "1111100010110011",
    "1111100000001010",
    "1111011101001100",
    "1111011010001001",
    "1111010111010000",
    "1111010100101010",
    "1111010010011100",
    "1111010000011110",
    "1111001110110001",
    "1111001101010110",
    "1111001100001111",
    "1111001011101010",
    "1111001011110010",
    "1111001100110111",
    "1111001110111111",
    "1111010010000101",
    "1111010101111110",
    "1111011010011000",
    "1111011110111111",
    "1111100011011111",
    "1111100111101110",
    "1111101011100100",
    "1111101110111101",
    "1111110001111100",
    "1111110100100010",
    "1111110110110001",
    "1111111000101101",
    "1111111010010110",
    "1111111011110000",
    "1111111101000101",
    "1111111110100100",
    "1111111111011011",
    "1111111100100000",
    "1111111000001011",
    "1111110010000110",
    "1111101010000100",
    "1111100000010001",
    "1111010101001001",
    "1111001001100101",
    "1110111110011100",
    "1110110100101111",
    "1110101101001001",
    "1110100111111100",
    "1110100101000110",
    "1110100100010000",
    "1110100100110111",
    "1110100110011111",
    "1110101000101101",
    "1110101011010110",
    "1110101110010110",
    "1110110001101011",
    "1110110101010010",
    "1110111001000110",
    "1110111101000000",
    "1111000000110110",
    "1111000100011100",
    "1111000111100010",
    "1111001001111111",
    "1111001011100011",
    "1111001100000010",
    "1111001011010100",
    "1111001001011110",
    "1111000110101100",
    "1111000011010010",
    "1110111111101001",
    "1110111100001110",
    "1110111001010001",
    "1110110111000011",
    "1110110101100100",
    "1110110100110110",
    "1110110100110100",
    "1110110101011000",
    "1110110110011011",
    "1110110111111111",
    "1110111010000010",
    "1110111100100110",
    "1110111111101011",
    "1111000011010010",
    "1111000111011000",
    "1111001011111100",
    "1111010000111011",
    "1111010110010011",
    "1111011100001010",
    "1111100010100111",
    "1111101001111000",
    "1111110010001100",
    "1111111011101101",
    "1111111001100110",
    "1111101110000110",
    "1111100010011001",
    "1111010111010000",
    "1111001101010100",
    "1111000101000001",
    "1110111110011001",
    "1110111001000111",
    "1110110100101100",
    "1110110000100100",
    "1110101100011001",
    "1110101000000011",
    "1110100011100110",
    "1110011111010010",
    "1110011011011101",
    "1110011000010101",
    "1110010110001110",
    "1110010101010101",
    "1110010101110010",
    "1110010111101000",
    "1110011010110101",
    "1110011111010010",
    "1110100100111011",
    "1110101011100101",
    "1110110011000011",
    "1110111011001010",
    "1111000011101001",
    "1111001100001010",
    "1111010100011000",
    "1111011011110111",
    "1111100010001011",
    "1111100110111110",
    "1111101010001000",
    "1111101011101100",
    "1111101011110110",
    "1111101010111101",
    "1111101001011001",
    "1111100111100000",
    "1111100101011111",
    "1111100011011111",
    "1111100001100100",
    "1111011111110001",
    "1111011110010001",
    "1111011101000100",
    "1111011100010111",
    "1111011100010011",
    "1111011100111010",
    "1111011110001100",
    "1111100000000101",
    "1111100010100001",
    "1111100101010111",
    "1111101000100001",
    "1111101011111010",
    "1111101111100000",
    "1111110011001010",
    "1111110110110011",
    "1111111010010110",
    "1111111101101011",
    "1111111111010111",
    "1111111100111101",
    "1111111011010001",
    "1111111010011001",
    "1111111010011001",
    "1111111011010011",
    "1111111101000100",
    "1111111111101010",
    "1111111100111010",
    "1111111000101101",
    "1111110011101100",
    "1111101101110100",
    "1111100110111111",
    "1111011111001111",
    "1111010110100000",
    "1111001101000000",
    "1111000011000110",
    "1110111001010001",
    "1110110000001000",
    "1110101000010001",
    "1110100010000110",
    "1110011101110010",
    "1110011011010011",
    "1110011010011011",
    "1110011010111010",
    "1110011100100001",
    "1110011111000100",
    "1110100010100010",
    "1110100110111011",
    "1110101100001100",
    "1110110010010100",
    "1110111001001001",
    "1111000000100001",
    "1111001000001011",
    "1111001111111010",
    "1111010111011011",
    "1111011110011110",
    "1111100100110111",
    "1111101010011010",
    "1111101110111100",
    "1111110010011101",
    "1111110101000010",
    "1111110110110111",
    "1111111000000110",
    "1111111000110111",
    "1111111001001100",
    "1111111000111111",
    "1111111000000110",
    "1111110110010111",
    "1111110011101000",
    "1111101111110101",
    "1111101010111101",
    "1111100101000101",
    "1111011110011011",
    "1111010111010011",
    "1111010000001111",
    "1111001001111001",
    "1111000100110001",
    "1111000001010100",
    "1110111111100110",
    "1110111111011110",
    "1111000000100100",
    "1111000010100110",
    "1111000101010111",
    "1111001000110101",
    "1111001101010001",
    "1111010010110001",
    "1111011001011110",
    "1111100001010100",
    "1111101001111100",
    "1111110011000000",
    "1111111100000011",
    "1111111011010110",
    "1111110011100100",
    "1111101100110010",
    "1111100111001100",
    "1111100010111001",
    "1111100000000011",
    "1111011110110001",
    "1111011111001101",
    "1111100001100001",
    "1111100101101111",
    "1111101011111111",
    "1111110100001010",
    "1111111110000011",
    "1111110110110000",
    "1111101011000011",
    "1111011111101100",
    "1111010101101001",
    "1111001101100011",
    "1111000111110111",
    "1111000100011101",
    "1111000010111110",
    "1111000010110001",
    "1111000011010000",
    "1111000100000011",
    "1111000101000101",
    "1111000110011111",
    "1111001000100010",
    "1111001011011101",
    "1111001111001111",
    "1111010011110001",
    "1111011000101101",
    "1111011101101110",
    "1111100010100100",
    "1111100110111110",
    "1111101010111100",
    "1111101110011101",
    "1111110001100110",
    "1111110100011100",
    "1111110111000101",
    "1111111001101001",
    "1111111100001101",
    "1111111110110110",
    "1111111110010001",
    "1111111011001101",
    "1111110111111010",
    "1111110100011000",
    "1111110000110011",
    "1111101101011000",
    "1111101010011110",
    "1111101000011101",
    "1111100111101101",
    "1111101000011011",
    "1111101010100111",
    "1111101110000111",
    "1111110010100011",
    "1111110111100101",
    "1111111100111010",
    "1111111101101011",
    "1111111000011010",
    "1111110011011010",
    "1111101110111011",
    "1111101011010000",
    "1111101000101011",
    "1111100111011001",
    "1111100111100010",
    "1111101000111111",
    "1111101011100100",
    "1111101111000100",
    "1111110011010010",
    "1111111000000111",
    "1111111101011100",
    "1111111100101111",
    "1111110110101000",
    "1111110000010100",
    "1111101010000000",
    "1111100011110110",
    "1111011110000100",
    "1111011000110010",
    "1111010100001000",
    "1111010000001100",
    "1111001101000100",
    "1111001010110010",
    "1111001001011011",
    "1111001000111010",
    "1111001001001100",
    "1111001010001011",
    "1111001011101010",
    "1111001101100000",
    "1111001111011100",
    "1111010001010100",
    "1111010010110100",
    "1111010011101110",
    "1111010011100100",
    "1111010010000000",
    "1111001110100100",
    "1111001001000010",
    "1111000001011010",
    "1110111000000001",
    "1110101101100001",
    "1110100010101111",
    "1110011000100010",
    "1110001111100011",
    "1110001000001100",
    "1110000010100111",
    "1101111110101001",
    "1101111011111111",
    "1101111010011000",
    "1101111001011011",
    "1101111000111111",
    "1101111000111010",
    "1101111001000110",
    "1101111001100111",
    "1101111010011110",
    "1101111011111100",
    "1101111110000111",
    "1110000001010101",
    "1110000101110100",
    "1110001011101011",
    "1110010011000000",
    "1110011011100001",
    "1110100100110111",
    "1110101110011100",
    "1110110111101100",
    "1111000000001101",
    "1111000111110101",
    "1111001110110001",
    "1111010101011000",
    "1111011100000111",
    "1111100011010010",
    "1111101010111110",
    "1111110011000001",
    "1111111011000100",
    "1111111101010001",
    "1111110110011011",
    "1111110000101001",
    "1111101011111110",
    "1111101000011001",
    "1111100101110001",
    "1111100011111001",
    "1111100010101100",
    "1111100010000011",
    "1111100001111101",
    "1111100010010111",
    "1111100011010101",
    "1111100100111001",
    "1111100111000100",
    "1111101001111000",
    "1111101101010010",
    "1111110001001100",
    "1111110101011001",
    "1111111001100101",
    "1111111101011110",
    "1111111111001111",
    "1111111100111010",
    "1111111011101010",
    "1111111011100011",
    "1111111100011110",
    "1111111110001110",
    "1111111111011001",
    "1111111100110000",
    "1111111001111111",
    "1111110111010101",
    "1111110100110110",
    "1111110010101101",
    "1111110000111110",
    "1111101111101100",
    "1111101110111011",
    "1111101110101000",
    "1111101110101111",
    "1111101111001100",
    "1111110000000000",
    "1111110001010000",
    "1111110011000001",
    "1111110101011011",
    "1111111000100010",
    "1111111100010100",
    "1111111111010110",
    "1111111010110010",
    "1111110110001110",
    "1111110010000000",
    "1111101110011001",
    "1111101011100100",
    "1111101001101000",
    "1111101000100011",
    "1111101000001110",
    "1111101000011011",
    "1111101000111100",
    "1111101001100100",
    "1111101010001101",
    "1111101010110111",
    "1111101011101001",
    "1111101100100110",
    "1111101101101110",
    "1111101110111011",
    "1111101111111110",
    "1111110000100011",
    "1111110000011001",
    "1111101111001111",
    "1111101100111110",
    "1111101001100010",
    "1111100101000101",
    "1111011111101110",
    "1111011001110000",
    "1111010011011100",
    "1111001101000000",
    "1111000110101100",
    "1111000000100110",
    "1110111010110101",
    "1110110101011111",
    "1110110000100110",
    "1110101100010100",
    "1110101000101101",
    "1110100101111100",
    "1110100100000110",
    "1110100011001010",
    "1110100011000101",
    "1110100011101100",
    "1110100100110100",
    "1110100110010110",
    "1110101000001011",
    "1110101010001100",
    "1110101100011110",
    "1110101110111011",
    "1110110001100010",
    "1110110100001110",
    "1110110110111001",
    "1110111001011101",
    "1110111011111100",
    "1110111110010111",
    "1111000000111000",
    "1111000011101100",
    "1111000110111011",
    "1111001010101011",
    "1111001111000100",
    "1111010100000000",
    "1111011001011011",
    "1111011111001101",
    "1111100101010000",
    "1111101011011000",
    "1111110001011001",
    "1111110111000101",
    "1111111100001110",
    "1111111111010100",
    "1111111011101111",
    "1111111000111111",
    "1111110110111101",
    "1111110101011110",
    "1111110100010011",
    "1111110011001100",
    "1111110001111111",
    "1111110000100011",
    "1111101110110110",
    "1111101100111001",
    "1111101010101101",
    "1111101000010110",
    "1111100101110010",
    "1111100011000000",
    "1111011111110110",
    "1111011100010001",
    "1111011000001011",
    "1111010011101010",
    "1111001110111011",
    "1111001010001100",
    "1111000101110001",
    "1111000001110011",
    "1110111110010010",
    "1110111011001110",
    "1110111000011011",
    "1110110101110110",
    "1110110011100010",
    "1110110001110001",
    "1110110000110000",
    "1110110000101110",
    "1110110001101110",
    "1110110011101001",
    "1110110110001110",
    "1110111001000110",
    "1110111011110101",
    "1110111110000111",
    "1110111111110000",
    "1111000000100111",
    "1111000000110011",
    "1111000000011001",
    "1110111111100100",
    "1110111110011011",
    "1110111101000000",
    "1110111011011001",
    "1110111001100101",
    "1110110111100111",
    "1110110101101001",
    "1110110011111100",
    "1110110010110001",
    "1110110010010101",
    "1110110010110011",
    "1110110100000001",
    "1110110101111011",
    "1110111000001011",
    "1110111010100011",
    "1110111100111000",
    "1110111111000111",
    "1111000001010000",
    "1111000011011000",
    "1111000101100101",
    "1111000111111001",
    "1111001010001100",
    "1111001100011001",
    "1111001110010001",
    "1111001111101000",
    "1111010000010100",
    "1111010000001101",
    "1111001111011001",
    "1111001101110111",
    "1111001011101010",
    "1111001000110111",
    "1111000101100010",
    "1111000001110001",
    "1110111101110011",
    "1110111010000001",
    "1110110110110110",
    "1110110100101110",
    "1110110011111011",
    "1110110100100010",
    "1110110110011010",
    "1110111001010000",
    "1110111100101010",
    "1111000000010010",
    "1111000011110100",
    "1111000111000011",
    "1111001001101101",
    "1111001011101000",
    "1111001100100110",
    "1111001100100000",
    "1111001011010100",
    "1111001001001011",
    "1111000110010000",
    "1111000010111000",
    "1110111111010100",
    "1110111011111000",
    "1110111000110101",
    "1110110110011011",
    "1110110100111110",
    "1110110100101111",
    "1110110110000000",
    "1110111000111111",
    "1110111101110101",
    "1111000100011111",
    "1111001100101000",
    "1111010101110001",
    "1111011111001010",
    "1111101000000011",
    "1111101111101100",
    "1111110101100110",
    "1111111001100011",
    "1111111011101000",
    "1111111100000100",
    "1111111011001101",
    "1111111001010100",
    "1111110110100100",
    "1111110011000001",
    "1111101110101111",
    "1111101001110100",
    "1111100100011111",
    "1111011111000111",
    "1111011010000111",
    "1111010110000001",
    "1111010011001010",
    "1111010001110001",
    "1111010001111011",
    "1111010011100111",
    "1111010110101111",
    "1111011011001010",
    "1111100000110001",
    "1111100111010100",
    "1111101110011100",
    "1111110101100111",
    "1111111100001000",
    "1111111110101100",
    "1111111011100010",
    "1111111010101001",
    "1111111011111110",
    "1111111111001100",
    "1111111100001011",
    "1111110110110111",
    "1111110001011100",
    "1111101100011001",
    "1111101000001010",
    "1111100100111011",
    "1111100010101110",
    "1111100001011001",
    "1111100000101011",
    "1111100000010010",
    "1111011111111111",
    "1111011111101001",
    "1111011111001101",
    "1111011110110000",
    "1111011110011100",
    "1111011110010111",
    "1111011110101001",
    "1111011111010111",
    "1111100000011110",
    "1111100001111011",
    "1111100011101110",
    "1111100101110001",
    "1111101000000100",
    "1111101010100101",
    "1111101101010100",
    "1111110000010000",
    "1111110011011011",
    "1111110110110111",
    "1111111010101100",
    "1111111110111110",
    "1111111100001010",
    "1111110110110001",
    "1111110000111010",
    "1111101010110001",
    "1111100100101001",
    "1111011110110110",
    "1111011001110000",
    "1111010101100101",
    "1111010010010111",
    "1111010000000011",
    "1111001110010111",
    "1111001101000100",
    "1111001011110011",
    "1111001010010001",
    "1111001000010011",
    "1111000101110110",
    "1111000010110110",
    "1110111111011110",
    "1110111011110111",
    "1110111000010000",
    "1110110100111100",
    "1110110010010100",
    "1110110000101110",
    "1110110000101001",
    "1110110010011010",
    "1110110110001110",
    "1110111100001010",
    "1111000100000110",
    "1111001101110010",
    "1111011000101101",
    "1111100100010010",
    "1111101111101010",
    "1111111001111010",
    "1111111101110000",
    "1111110111111110",
    "1111110100110111",
    "1111110100001111",
    "1111110101100101",
    "1111111000010001",
    "1111111011110000",
    "1111111111101010",
    "1111111100001001",
    "1111110111110001",
    "1111110011001101",
    "1111101110100001",
    "1111101001110011",
    "1111100101001110",
    "1111100000111000",
    "1111011100110011",
    "1111011000111010",
    "1111010101000000",
    "1111010000110011",
    "1111001100000001",
    "1111000110011011",
    "1111000000000101",
    "1110111001001001",
    "1110110010000101",
    "1110101011011000",
    "1110100101011101",
    "1110100000100100",
    "1110011100110010",
    "1110011001111010",
    "1110010111101111",
    "1110010110001001",
    "1110010101001000",
    "1110010100101010",
    "1110010100110110",
    "1110010101100100",
    "1110010110101100",
    "1110010111111100",
    "1110011001001100",
    "1110011010010011",
    "1110011011011000",
    "1110011100100011",
    "1110011110001001",
    "1110100000010100",
    "1110100011010000",
    "1110100110111110",
    "1110101011001111",
    "1110101111110101",
    "1110110100011000",
    "1110111000100101",
    "1110111100001111",
    "1110111111001111",
    "1111000001100100",
    "1111000011010111",
    "1111000100101110",
    "1111000101111001",
    "1111000110111111",
    "1111001000001011",
    "1111001001100011",
    "1111001011001110",
    "1111001101010010",
    "1111001111111010",
    "1111010011001011",
    "1111010111001110",
    "1111011011111101",
    "1111100001010101",
    "1111100111000111",
    "1111101100111111",
    "1111110010101011",
    "1111110111111100",
    "1111111100101001",
    "1111111111001010",
    "1111111011011100",
    "1111110111111100",
    "1111110100011111",
    "1111110000111010",
    "1111101101001101",
    "1111101001011100",
    "1111100101110110",
    "1111100010101011",
    "1111100000001100",
    "1111011110100011",
    "1111011101110101",
    "1111011101111000",
    "1111011110100001",
    "1111011111011110",
    "1111100000010111",
    "1111100001000000",
    "1111100001001111",
    "1111100000111101",
    "1111100000001100",
    "1111011110111111",
    "1111011101011100",
    "1111011011101010",
    "1111011001101111",
    "1111010111101101",
    "1111010101101010",
    "1111010011100110",
    "1111010001100110",
    "1111001111101001",
    "1111001101111000",
    "1111001100010011",
    "1111001010111100",
    "1111001001110101",
    "1111001000111110",
    "1111001000011011",
    "1111001000010011",
    "1111001000110010",
    "1111001010000110",
    "1111001100010110",
    "1111001111101001",
    "1111010011110011",
    "1111011000011110",
    "1111011101001100",
    "1111100001010111",
    "1111100100011111",
    "1111100110001110",
    "1111100110100111",
    "1111100101110111",
    "1111100100011101",
    "1111100010111110",
    "1111100001111000",
    "1111100001100110",
    "1111100010010101",
    "1111100100010000",
    "1111100111011001",
    "1111101011110100",
    "1111110001100110",
    "1111111000111001",
    "1111111110000110",
    "1111110011011001",
    "1111100111001001",
    "1111011001111100",
    "1111001100101110",
    "1111000000100100",
    "1110110110011111",
    "1110101111000101",
    "1110101010011110",
    "1110101000010101",
    "1110100111111111",
    "1110101000110111",
    "1110101010100010",
    "1110101100110010",
    "1110101111110011",
    "1110110011101100",
    "1110111000100101",
    "1110111110010111",
    "1111000100101100",
    "1111001010111101",
    "1111010000100011",
    "1111010100101100",
    "1111010110110110",
    "1111010110101100",
    "1111010100001011",
    "1111001111101000",
    "1111001001101000",
    "1111000011000001",
    "1110111100101000",
    "1110110111001000",
    "1110110010111000",
    "1110110000000000",
    "1110101110010110",
    "1110101101100110",
    "1110101101011110",
    "1110101101101011",
    "1110101110000111",
    "1110101110101001",
    "1110101111010010",
    "1110110000000111",
    "1110110001001100",
    "1110110010101001",
    "1110110100101001",
    "1110110111010101",
    "1110111010110000",
    "1110111110111010",
    "1111000011101010",
    "1111001000110101",
    "1111001110010111",
    "1111010100001000",
    "1111011010001111",
    "1111100000111011",
    "1111101000010101",
    "1111110000101001",
    "1111111001111100",
    "1111111011110010",
    "1111110000110111",
    "1111100101100100",
    "1111011010011001",
    "1111001111111011",
    "1111000110100101",
    "1110111110101110",
    "1110111000011110",
    "1110110011101111",
    "1110110000001111",
    "1110101101100000",
    "1110101011000111",
    "1110101000101111",
    "1110100110001011",
    "1110100011011101",
    "1110100000110001",
    "1110011110011011",
    "1110011100110101",
    "1110011100011011",
    "1110011101011110",
    "1110100000001000",
    "1110100100011010",
    "1110101010000111",
    "1110110001000011",
    "1110111000111111",
    "1111000001100110",
    "1111001010101000",
    "1111010011101010",
    "1111011100001100",
    "1111100011100100",
    "1111101001001110",
    "1111101100110101",
    "1111101110011011",
    "1111101110011001",
    "1111101101011000",
    "1111101100000100",
    "1111101011000000",
    "1111101010011011",
    "1111101010010001",
    "1111101010010011",
    "1111101010001110",
    "1111101001111000",
    "1111101001010010",
    "1111101000101100",
    "1111101000011100",
    "1111101000111000",
    "1111101010001101",
    "1111101100011110",
    "1111101111100100",
    "1111110011010011",
    "1111110111011101",
    "1111111011110010",
    "1111111111110111",
    "1111111011110001",
    "1111111000000101",
    "1111110100111101",
    "1111110010100100",
    "1111110001000010",
    "1111110000011011",
    "1111110000110001",
    "1111110010000010",
    "1111110100001010",
    "1111110111000011",
    "1111111010101100",
    "1111111111000000",
    "1111111011111100",
    "1111110110001101",
    "1111101111101011",
    "1111101000001111",
    "1111011111110011",
    "1111010110010101",
    "1111001100000001",
    "1111000001001111",
    "1110110110101101",
    "1110101101001111",
    "1110100101100100",
    "1110100000001000",
    "1110011101000111",
    "1110011100001111",
    "1110011101000010",
    "1110011110111101",
    "1110100001100100",
    "1110100100101001",
    "1110101000001011",
    "1110101100011011",
    "1110110001100010",
    "1110110111101101",
    "1110111110111000",
    "1111000110110100",
    "1111001111001010",
    "1111010111011011",
    "1111011111000111",
    "1111100101110100",
    "1111101011010010",
    "1111101111011011",
    "1111110010010110",
    "1111110100010000",
    "1111110101011010",
    "1111110101111111",
    "1111110110000100",
    "1111110101101000",
    "1111110100100010",
    "1111110010100110",
    "1111101111101001",
    "1111101011011110",
    "1111100101111110",
    "1111011111001000",
    "1111010111001011",
    "1111001110100011",
    "1111000101111001",
    "1110111101111101",
    "1110110111011000",
    "1110110010100111",
    "1110101111110101",
    "1110101110110110",
    "1110101111100001",
    "1110110001011111",
    "1110110100100111",
    "1110111000110100",
    "1110111110001001",
    "1111000100100100",
    "1111001100000010",
    "1111010100010011",
    "1111011100111101",
    "1111100101100010",
    "1111101101101000",
    "1111110100111110",
    "1111111011011111",
    "1111111110101111",
    "1111111001101100",
    "1111110101010010",
    "1111110001100011",
    "1111101110101000",
    "1111101100110010",
    "1111101100001111",
    "1111101101001111",
    "1111101111111000",
    "1111110100010011",
    "1111111010100001",
    "1111111101100001",
    "1111110100001010",
    "1111101001111001",
    "1111011111100011",
    "1111010101111100",
    "1111001101111000",
    "1111000111110001",
    "1111000011101010",
    "1111000001010000",
    "1111000000000101",
    "1110111111101001",
    "1110111111101011",
    "1111000000000011",
    "1111000000111011",
    "1111000010011101",
    "1111000100110001",
    "1111000111111010",
    "1111001011110000",
    "1111010000000011",
    "1111010100100000",
    "1111011000110111",
    "1111011100111000",
    "1111100000011010",
    "1111100011011100",
    "1111100101111100",
    "1111101000000111",
    "1111101010000111",
    "1111101100001111",
    "1111101110101110",
    "1111110001101101",
    "1111110101010100",
    "1111111001100101",
    "1111111110011100",
    "1111111100000100",
    "1111110110000011",
    "1111101111100100",
    "1111101000111001",
    "1111100010011100",
    "1111011100111010",
    "1111011001000010",
    "1111010111101000",
    "1111011001010001",
    "1111011110001100",
    "1111100110001001",
    "1111110000011111",
    "1111111100000111",
    "1111111000001111",
    "1111101101111001",
    "1111100101110100",
    "1111100000100110",
    "1111011110010010",
    "1111011110100001",
    "1111100000101011",
    "1111100100000000",
    "1111100111111111",
    "1111101100010100",
    "1111110000111000",
    "1111110101110010",
    "1111111011001001",
    "1111111110111100",
    "1111111000100110",
    "1111110010000000",
    "1111101011011111",
    "1111100101011010",
    "1111100000000010",
    "1111011011100011",
    "1111011000000001",
    "1111010101011010",
    "1111010011101001",
    "1111010010100110",
    "1111010010010000",
    "1111010010100010",
    "1111010011011010",
    "1111010100101110",
    "1111010110001001",
    "1111010111011011",
    "1111011000010000",
    "1111011000011000",
    "1111010111101101",
    "1111010110010000",
    "1111010100000101",
    "1111010001001111",
    "1111001101101101",
    "1111001001011000",
    "1111000100001011",
    "1110111101111101",
    "1110110110101111",
    "1110101110100110",
    "1110100101110001",
    "1110011100101101",
    "1110010011110110",
    "1110001011110011",
    "1110000101000000",
    "1101111111110011",
    "1101111100010110",
    "1101111010100011",
    "1101111010001100",
    "1101111010111111",
    "1101111100100011",
    "1101111110100110",
    "1110000000110011",
    "1110000010111110",
    "1110000100111011",
    "1110000110101100",
    "1110001000011000",
    "1110001010001111",
    "1110001100101010",
    "1110010000000010",
    "1110010100100111",
    "1110011010100011",
    "1110100001101110",
    "1110101001110010",
    "1110110010010000",
    "1110111010101010",
    "1111000010101001",
    "1111001010000001",
    "1111010000110011",
    "1111010111001101",
    "1111011101011100",
    "1111100011110001",
    "1111101010001110",
    "1111110000101111",
    "1111110111000101",
    "1111111100111100",
    "1111111110000000",
    "1111111010000010",
    "1111110111010100",
    "1111110101110100",
    "1111110101011001",
    "1111110101110011",
    "1111110110101111",
    "1111110111111000",
    "1111111001000000",
    "1111111001111000",
    "1111111010011100",
    "1111111010101110",
    "1111111010110110",
    "1111111010111111",
    "1111111011010000",
    "1111111011110000",
    "1111111100011111",
    "1111111101010101",
    "1111111110001100",
    "1111111110111010",
    "1111111111011001",
    "1111111111100101",
    "1111111111011110",
    "1111111110111110",
    "1111111110000100",
    "1111111100101100",
    "1111111010110111",
    "1111111000101001",
    "1111110110001100",
    "1111110011101101",
    "1111110001011010",
    "1111101111100010",
    "1111101110001110",
    "1111101101101000",
    "1111101101110100",
    "1111101110110001",
    "1111110000100000",
    "1111110010111010",
    "1111110101111001",
    "1111111001010100",
    "1111111101000001",
    "1111111111000011",
    "1111111011000011",
    "1111110111000000",
    "1111110010111110",
    "1111101111000011",
    "1111101011011010",
    "1111101000010010",
    "1111100101111001",
    "1111100100011101",
    "1111100100001011",
    "1111100101000001",
    "1111100110110111",
    "1111101001011100",
    "1111101100011001",
    "1111101111010111",
    "1111110001111111",
    "1111110100000011",
    "1111110101011000",
    "1111110101111000",
    "1111110101100000",
    "1111110100001110",
    "1111110010000110",
    "1111101111001100",
    "1111101011101101",
    "1111100111110110",
    "1111100011111001",
    "1111011111111111",
    "1111011100010011",
    "1111011000110010",
    "1111010101011000",
    "1111010001111011",
    "1111001110010010",
    "1111001010011001",
    "1111000110010101",
    "1111000010001111",
    "1110111110010001",
    "1110111010101010",
    "1110110111100010",
    "1110110100111110",
    "1110110011000000",
    "1110110001100100",
    "1110110000101001",
    "1110110000001010",
    "1110110000001000",
    "1110110000100100",
    "1110110001011010",
    "1110110010101110",
    "1110110100011100",
    "1110110110011101",
    "1110111000101101",
    "1110111011000110",
    "1110111101100011",
    "1111000000000010",
    "1111000010100010",
    "1111000101001011",
    "1111001000000100",
    "1111001011010100",
    "1111001111000101",
    "1111010011011111",
    "1111011000100011",
    "1111011110010100",
    "1111100100101001",
    "1111101011010011",
    "1111110010000011",
    "1111111000100101",
    "1111111110100111",
    "1111111100000011",
    "1111110111101000",
    "1111110100001101",
    "1111110001110110",
    "1111110000100100",
    "1111110000010010",
    "1111110000110111",
    "1111110010000010",
    "1111110011011101",
    "1111110100101110",
    "1111110101100000",
    "1111110101011101",
    "1111110100010111",
    "1111110010000110",
    "1111101110101010",
    "1111101010000111",
    "1111100100101001",
    "1111011110011100",
    "1111010111110100",
    "1111010001000101",
    "1111001010100101",
    "1111000100100101",
    "1110111111010110",
    "1110111011000100",
    "1110110111111010",
    "1110110101111100",
    "1110110101001101",
    "1110110101100111",
    "1110110111001001",
    "1110111001100101",
    "1110111100110010",
    "1111000000011001",
    "1111000100000011",
    "1111000111010110",
    "1111001001110111",
    "1111001011010001",
    "1111001011011001",
    "1111001010010011",
    "1111001000001000",
    "1111000101001101",
    "1111000001110000",
    "1110111101111101",
    "1110111001111010",
    "1110110101101100",
    "1110110001011001",
    "1110101101001111",
    "1110101001100011",
    "1110100110101111",
    "1110100101001101",
    "1110100101001110",
    "1110100110111011",
    "1110101010001011",
    "1110101110101110",
    "1110110100001011",
    "1110111010000111",
    "1111000000000111",
    "1111000101101110",
    "1111001010101010",
    "1111001110101011",
    "1111010001101011",
    "1111010011101010",
    "1111010100110001",
    "1111010101001001",
    "1111010101000000",
    "1111010100100000",
    "1111010011110110",
    "1111010011000101",
    "1111010010001101",
    "1111010001001101",
    "1111001111111010",
    "1111001110001100",
    "1111001011111100",
    "1111001001001011",
    "1111000110001000",
    "1111000011001000",
    "1111000000101100",
    "1110111111001111",
    "1110111111000010",
    "1111000000001010",
    "1111000010100001",
    "1111000101110001",
    "1111001001100000",
    "1111001101010110",
    "1111010000110110",
    "1111010011101010",
    "1111010101011010",
    "1111010101110100",
    "1111010100100101",
    "1111010001101001",
    "1111001101001001",
    "1111000111011101",
    "1111000001001111",
    "1110111011001001",
    "1110110101111110",
    "1110110010001111",
    "1110110000001101",
    "1110101111111010",
    "1110110001000011",
    "1110110011010101",
    "1110110110011101",
    "1110111010010011",
    "1110111110110110",
    "1111000100001110",
    "1111001010100000",
    "1111010001100111",
    "1111011001010101",
    "1111100001000101",
    "1111101000010100",
    "1111101110011001",
    "1111110010110111",
    "1111110101011101",
    "1111110110001110",
    "1111110101011010",
    "1111110011011010",
    "1111110000101111",
    "1111101101111101",
    "1111101011011111",
    "1111101001101110",
    "1111101000110101",
    "1111101000111001",
    "1111101001110101",
    "1111101011100001",
    "1111101101110000",
    "1111110000010111",
    "1111110011001010",
    "1111110110000010",
    "1111111000111000",
    "1111111011100110",
    "1111111110001100",
    "1111111111011000",
    "1111111101001111",
    "1111111011011010",
    "1111111010000000",
    "1111111001000100",
    "1111111000101000",
    "1111111000101101",
    "1111111001010000",
    "1111111010010011",
    "1111111011110111",
    "1111111110000000",
    "1111111111001001",
    "1111111011100100",
    "1111110111001111",
    "1111110010010101",
    "1111101101001000",
    "1111100111111111",
    "1111100011010000",
    "1111011111001000",
    "1111011011101101",
    "1111011000111010",
    "1111010110100101",
    "1111010100100000",
    "1111010010100010",
    "1111010000101100",
    "1111001111000111",
    "1111001101111111",
    "1111001101100110",
    "1111001110001111",
    "1111001111111111",
    "1111010010110011",
    "1111010110100010",
    "1111011010111100",
    "1111011111101001",
    "1111100100011100",
    "1111101000111111",
    "1111101101001011",
    "1111110000111110",
    "1111110100011101",
    "1111110111110111",
    "1111111011011101",
    "1111111111100010",
    "1111111011100110",
    "1111110101110110",
    "1111101111010000",
    "1111101000000011",
    "1111100000101001",
    "1111011001100000",
    "1111010011000110",
    "1111001101110010",
    "1111001001101111",
    "1111000110111111",
    "1111000101100100",
    "1111000101010000",
    "1111000101110111",
    "1111000111001001",
    "1111001000110000",
    "1111001010011000",
    "1111001011110010",
    "1111001100110000",
    "1111001101010100",
    "1111001101100011",
    "1111001101101101",
    "1111001110000000",
    "1111001110111010",
    "1111010000101100",
    "1111010011101111",
    "1111011000010110",
    "1111011110100100",
    "1111100110010101",
    "1111101111001101",
    "1111111000100100",
    "1111111110010101",
    "1111110110011000",
    "1111110000000111",
    "1111101011110110",
    "1111101001100111",
    "1111101001001011",
    "1111101010001100",
    "1111101100010101",
    "1111101111010010",
    "1111110010111010",
    "1111110111000101",
    "1111111011101101",
    "1111111111010011",
    "1111111010001110",
    "1111110101001101",
    "1111110000011110",
    "1111101100001111",
    "1111101000100100",
    "1111100101011010",
    "1111100010101011",
    "1111100000000111",
    "1111011101011110",
    "1111011010100000",
    "1111010110110111",
    "1111010010010101",
    "1111001100101101",
    "1111000101111001",
    "1110111110000010",
    "1110110101100010",
    "1110101100111100",
    "1110100100110111",
    "1110011101111011",
    "1110011000100111",
    "1110010101000011",
    "1110010011001111",
    "1110010010111011",
    "1110010011110001",
    "1110010101011011",
    "1110010111101100",
    "1110011010010110",
    "1110011101011001",
    "1110100000110001",
    "1110100100011101",
    "1110101000010000",
    "1110101011111111",
    "1110101111011001",
    "1110110010001011",
    "1110110100001110",
    "1110110101100000",
    "1110110110001000",
    "1110110110010010",
    "1110110110001011",
    "1110110110000011",
    "1110110110000001",
    "1110110110001011",
    "1110110110100010",
    "1110110111000100",
    "1110110111110111",
    "1110111001000010",
    "1110111010110101",
    "1110111101010111",
    "1111000000110110",
    "1111000101001101",
    "1111001010010011",
    "1111001111111101",
    "1111010101111011",
    "1111011011111111",
    "1111100010000010",
    "1111100111111111",
    "1111101101110100",
    "1111110011011101",
    "1111111000110010",
    "1111111101101010",
    "1111111110000010",
    "1111111010011001",
    "1111110111011000",
    "1111110100110100",
    "1111110010100110",
    "1111110000100110",
    "1111101110110100",
    "1111101101010110",
    "1111101100010011",
    "1111101011110001",
    "1111101011110000",
    "1111101100001001",
    "1111101100101011",
    "1111101101000110",
    "1111101101001000",
    "1111101100101010",
    "1111101011101011",
    "1111101010001111",
    "1111101000011100",
    "1111100110011101",
    "1111100100010010",
    "1111100001111110",
    "1111011111100001",
    "1111011100111101",
    "1111011010010110",
    "1111010111111010",
    "1111010101110100",
    "1111010100010000",
    "1111010011011100",
    "1111010011011101",
    "1111010100010011",
    "1111010101111100",
    "1111011000001011",
    "1111011010110101",
    "1111011101101011",
    "1111100000011010",
    "1111100010111000",
    "1111100100101111",
    "1111100101111001",
    "1111100110001001",
    "1111100101100000",
    "1111100100000110",
    "1111100010000011",
    "1111011111101011",
    "1111011101001111",
    "1111011011000010",
    "1111011001010011",
    "1111011000001110",
    "1111010111111100",
    "1111011000100111",
    "1111011010010110",
    "1111011101010110",
    "1111100001101110",
    "1111100111101000",
    "1111101111000101",
    "1111111000000100",
    "1111111101011010",
    "1111110001100011",
    "1111100100101100",
    "1111010111100000",
    "1111001010111111",
    "1111000000001101",
    "1110111000000011",
    "1110110010111101",
    "1110110000110000",
    "1110110000101110",
    "1110110001111000",
    "1110110011010010",
    "1110110100011000",
    "1110110101000000",
    "1110110101011000",
    "1110110101110111",
    "1110110110110010",
    "1110111000010110",
    "1110111010011101",
    "1110111100111000",
    "1110111111010110",
    "1111000001100010",
    "1111000011001011",
    "1111000100000000",
    "1111000011101100",
    "1111000010001000",
    "1110111111010001",
    "1110111011010011",
    "1110110110101010",
    "1110110001111000",
    "1110101101100100",
    "1110101010001001",
    "1110100111110111",
    "1110100110101101",
    "1110100110100010",
    "1110100110111111",
    "1110100111110100",
    "1110101000101111",
    "1110101001101010",
    "1110101010100101",
    "1110101011100110",
    "1110101100111101",
    "1110101110110101",
    "1110110001011110",
    "1110110100111110",
    "1110111001011101",
    "1110111110111011",
    "1111000101010010",
    "1111001100001111",
    "1111010011100001",
    "1111011010110100",
    "1111100001111000",
    "1111101000100110",
    "1111101111000010",
    "1111110101011000",
    "1111111011111101",
    "1111111100111001",
    "1111110100111111",
    "1111101100010100",
    "1111100011000001",
    "1111011001100000",
    "1111010000001111",
    "1111000111110001",
    "1111000000011110",
    "1110111010100101",
    "1110110110000110",
    "1110110010110100",
    "1110110000011100",
    "1110101110101000",
    "1110101101000111",
    "1110101011110011",
    "1110101010101000",
    "1110101001101011",
    "1110101001000100",
    "1110101000111001",
    "1110101001001100",
    "1110101010000111",
    "1110101011100101",
    "1110101101101101",
    "1110110000011100",
    "1110110011111000",
    "1110110111111110",
    "1110111100101110",
    "1111000010000110",
    "1111000111110111",
    "1111001101110011",
    "1111010011011010",
    "1111011000001100",
    "1111011011110000",
    "1111011101110011",
    "1111011110011011",
    "1111011101111000",
    "1111011100101000",
    "1111011011001110",
    "1111011001111111",
    "1111011001000110",
    "1111011000100111",
    "1111011000011011",
    "1111011000100010",
    "1111011000111111",
    "1111011001111111",
    "1111011011101011",
    "1111011110010010",
    "1111100001111110",
    "1111100110101110",
    "1111101100011001",
    "1111110010101110",
    "1111111001010110",
    "1111111111110100",
    "1111111010010001",
    "1111110101011011",
    "1111110001111100",
    "1111110000000000",
    "1111101111101110",
    "1111110000111111",
    "1111110011101001",
    "1111110111100001",
    "1111111100010111",
    "1111111101111111",
    "1111110111110010",
    "1111110001001010",
    "1111101010001111",
    "1111100011001010",
    "1111011011111100",
    "1111010100101100",
    "1111001101011110",
    "1111000110010011",
    "1110111111010111",
    "1110111000110010",
    "1110110010101111",
    "1110101101011001",
    "1110101000110010",
    "1110100101000000",
    "1110100010000000",
    "1110011111110000",
    "1110011110010001",
    "1110011101100100",
    "1110011101110000",
    "1110011110111000",
    "1110100001001000",
    "1110100100101111",
    "1110101001110101",
    "1110110000101011",
    "1110111001010011",
    "1111000011100010",
    "1111001110111010",
    "1111011010101011",
    "1111100101111011",
    "1111101111101100",
    "1111110111010000",
    "1111111100001111",
    "1111111110101011",
    "1111111110111011",
    "1111111101011111",
    "1111111010110110",
    "1111110111010110",
    "1111110011000010",
    "1111101101111001",
    "1111100111110011",
    "1111100000101011",
    "1111011000101010",
    "1111010000001101",
    "1111000111111010",
    "1111000000100001",
    "1110111010100101",
    "1110110110011101",
    "1110110100001011",
    "1110110011011000",
    "1110110011101010",
    "1110110100100000",
    "1110110101100111",
    "1110110110110110",
    "1110111000011000",
    "1110111010100011",
    "1110111101110010",
    "1111000010011100",
    "1111001000101101",
    "1111010000100100",
    "1111011001101011",
    "1111100011100001",
    "1111101101100000",
    "1111110111000111",
    "1111111111111101",
    "1111110111111111",
    "1111110001000000",
    "1111101011000100",
    "1111100110010011",
    "1111100010111011",
    "1111100001001101",
    "1111100001011010",
    "1111100011110001",
    "1111101000010000",
    "1111101110101100",
    "1111110110110000",
    "1111111111111000",
    "1111110110100001",
    "1111101101001100",
    "1111100100101111",
    "1111011101101011",
    "1111011000010000",
    "1111010100100000",
    "1111010010001101",
    "1111010001000000",
    "1111010000011100",
    "1111010000001111",
    "1111010000001101",
    "1111010000010010",
    "1111010000011111",
    "1111010000111001",
    "1111010001011111",
    "1111010010001101",
    "1111010011000000",
    "1111010011110100",
    "1111010100101010",
    "1111010101100111",
    "1111010110110010",
    "1111011000011010",
    "1111011010100011",
    "1111011101010001",
    "1111100000100011",
    "1111100100010011",
    "1111101000100001",
    "1111101101000110",
    "1111110010000010",
    "1111110111010100",
    "1111111100110110",
    "1111111101011010",
    "1111110111101011",
    "1111110010000111",
    "1111101100110111",
    "1111101000000111",
    "1111100011111100",
    "1111100000100110",
    "1111011110001111",
    "1111011101001010",
    "1111011101110010",
    "1111100000010100",
    "1111100101000110",
    "1111101100000100",
    "1111110100111011",
    "1111111110111000",
    "1111110111000111",
    "1111101110010110",
    "1111100111110101",
    "1111100100001101",
    "1111100011100110",
    "1111100101100100",
    "1111101001011001",
    "1111101110010100",
    "1111110011101011",
    "1111111001001011",
    "1111111110110000",
    "1111111011011011",
    "1111110101010101",
    "1111101110111101",
    "1111101000100010",
    "1111100010011010",
    "1111011101000000",
    "1111011000101100",
    "1111010101101001",
    "1111010011111011",
    "1111010011011111",
    "1111010100001011",
    "1111010101110110",
    "1111011000001110",
    "1111011011000110",
    "1111011110001010",
    "1111100001001010",
    "1111100011101110",
    "1111100101100111",
    "1111100110100010",
    "1111100110010101",
    "1111100100110110",
    "1111100010000101",
    "1111011110000111",
    "1111011001000100",
    "1111010011001011",
    "1111001100101000",
    "1111000101101100",
    "1110111110100110",
    "1110110111100000",
    "1110110000100111",
    "1110101010000010",
    "1110100011110011",
    "1110011101110011",
    "1110011000000011",
    "1110010010011001",
    "1110001100110101",
    "1110000111011101",
    "1110000010011010",
    "1101111101111010",
    "1101111010000110",
    "1101110111000100",
    "1101110100110111",
    "1101110011011010",
    "1101110010100110",
    "1101110010011001",
    "1101110010111000",
    "1101110100001110",
    "1101110110110010",
    "1101111010110101",
    "1110000000101100",
    "1110001000011101",
    "1110010010000000",
    "1110011101000100",
    "1110101001000110",
    "1110110101010101",
    "1111000001000010",
    "1111001011100000",
    "1111010100010101",
    "1111011011011001",
    "1111100000110101",
    "1111100101000101",
    "1111101000100110",
    "1111101011111000",
    "1111101111001110",
    "1111110010110100",
    "1111110110101010",
    "1111111010101101",
    "1111111110110101",
    "1111111101000010",
    "1111111001001010",
    "1111110101101100",
    "1111110010110001",
    "1111110000100101",
    "1111101111001110",
    "1111101110101110",
    "1111101110111111",
    "1111101111111000",
    "1111110001010000",
    "1111110010111101",
    "1111110100110101",
    "1111110110110001",
    "1111111000100111",
    "1111111010001110",
    "1111111011011001",
    "1111111011111101",
    "1111111011110010",
    "1111111010110011",
    "1111111001000001",
    "1111110110100010",
    "1111110011100100",
    "1111110000011001",
    "1111101101010011",
    "1111101010100100",
    "1111101000011001",
    "1111100110111010",
    "1111100110001001",
    "1111100110000100",
    "1111100110101000",
    "1111100111110000",
    "1111101001011000",
    "1111101011011111",
    "1111101110000000",
    "1111110000110111",
    "1111110011111010",
    "1111110111000000",
    "1111111001111100",
    "1111111100100101",
    "1111111110110101",
    "1111111111001111",
    "1111111101101000",
    "1111111100001010",
    "1111111010101010",
    "1111111001000011",
    "1111110111010110",
    "1111110101100110",
    "1111110100000011",
    "1111110010110110",
    "1111110010001011",
    "1111110010000110",
    "1111110010100011",
    "1111110011011001",
    "1111110100010110",
    "1111110101001101",
    "1111110101101111",
    "1111110101110110",
    "1111110101011101",
    "1111110100101010",
    "1111110011100001",
    "1111110010001100",
    "1111110000110000",
    "1111101111010000",
    "1111101101101010",
    "1111101011111000",
    "1111101001110011",
    "1111100111010111",
    "1111100100011101",
    "1111100001000111",
    "1111011101010110",
    "1111011001010000",
    "1111010100111011",
    "1111010000011110",
    "1111001100000001",
    "1111000111101000",
    "1111000011011101",
    "1110111111101000",
    "1110111100001010",
    "1110111001001110",
    "1110110110110001",
    "1110110100110011",
    "1110110011001101",
    "1110110001111011",
    "1110110000110110",
    "1110101111111111",
    "1110101111010010",
    "1110101110110101",
    "1110101110101101",
    "1110101110111111",
    "1110101111101100",
    "1110110000111011",
    "1110110010101011",
    "1110110101000000",
    "1110110111111001",
    "1110111011011000",
    "1110111111011111",
    "1111000100010010",
    "1111001001101101",
    "1111001111110000",
    "1111010110010010",
    "1111011101000000",
    "1111100011100111",
    "1111101001110001",
    "1111101111000100",
    "1111110011010001",
    "1111110110001111",
    "1111111000000010",
    "1111111000111000",
    "1111111001000001",
    "1111111000110100",
    "1111111000100111",
    "1111111000101000",
    "1111111001000101",
    "1111111010000110",
    "1111111011101101",
    "1111111110000010",
    "1111111110110100",
    "1111111010110110",
    "1111110110000001",
    "1111110000011001",
    "1111101010001000",
    "1111100011100001",
    "1111011100110010",
    "1111010110001101",
    "1111010000000000",
    "1111001010010011",
    "1111000101001000",
    "1111000000100100",
    "1110111100101101",
    "1110111001100111",
    "1110110111011011",
    "1110110110010110",
    "1110110110100100",
    "1110111000001001",
    "1110111011000100",
    "1110111111000111",
    "1111000011111011",
    "1111001000111010",
    "1111001101100011",
    "1111010001010000",
    "1111010011101110",
    "1111010100110100",
    "1111010100100100",
    "1111010011001011",
    "1111010000111001",
    "1111001101111111",
    "1111001010100011",
    "1111000110110001",
    "1111000010110001",
    "1110111110110101",
    "1110111011001110",
    "1110111000010110",
    "1110110110100100",
    "1110110110001001",
    "1110110111001101",
    "1110111001101011",
    "1110111101011011",
    "1111000010000010",
    "1111000111001001",
    "1111001100011011",
    "1111010001100001",
    "1111010110001000",
    "1111011010000010",
    "1111011101000100",
    "1111011111000111",
    "1111100000000011",
    "1111011111111010",
    "1111011110101011",
    "1111011100011011",
    "1111011001010101",
    "1111010101100000",
    "1111010001010010",
    "1111001100111010",
    "1111001000101111",
    "1111000101000101",
    "1111000010010100",
    "1111000000101001",
    "1111000000001101",
    "1111000000111110",
    "1111000010101110",
    "1111000101000110",
    "1111000111101000",
    "1111001001111001",
    "1111001011100011",
    "1111001100010111",
    "1111001100010111",
    "1111001011101010",
    "1111001010011001",
    "1111001000110111",
    "1111000111001110",
    "1111000101100101",
    "1111000100000000",
    "1111000010100100",
    "1111000001010101",
    "1111000000011100",
    "1111000000000000",
    "1111000000001010",
    "1111000001000011",
    "1111000010101100",
    "1111000100111100",
    "1111000111101100",
    "1111001010100011",
    "1111001101010001",
    "1111001111100011",
    "1111010001001111",
    "1111010010001101",
    "1111010010100001",
    "1111010010001111",
    "1111010001011110",
    "1111010000011100",
    "1111001111010111",
    "1111001110011110",
    "1111001110000000",
    "1111001110001111",
    "1111001111010001",
    "1111010001000111",
    "1111010011101010",
    "1111010110101100",
    "1111011001110100",
    "1111011100101010",
    "1111011110110110",
    "1111100000010001",
    "1111100000110110",
    "1111100000101100",
    "1111100000001000",
    "1111011111011111",
    "1111011111000100",
    "1111011111000111",
    "1111011111111000",
    "1111100001100001",
    "1111100100000110",
    "1111100111101011",
    "1111101100001010",
    "1111110001010100",
    "1111110110110001",
    "1111111100000101",
    "1111111111001101",
    "1111111011100101",
    "1111111001010010",
    "1111111000011011",
    "1111111001000010",
    "1111111011000100",
    "1111111110011010",
    "1111111101000000",
    "1111110111011110",
    "1111110001001111",
    "1111101010110010",
    "1111100100100100",
    "1111011111000100",
    "1111011010100010",
    "1111010111000100",
    "1111010100100111",
    "1111010010110110",
    "1111010001100100",
    "1111010000011111",
    "1111001111100011",
    "1111001110101000",
    "1111001101110010",
    "1111001100111111",
    "1111001100010100",
    "1111001011110010",
    "1111001011011000",
    "1111001011001010",
    "1111001011001010",
    "1111001011100000",
    "1111001100001111",
    "1111001101011110",
    "1111001111010100",
    "1111010001110100",
    "1111010101000001",
    "1111011000111111",
    "1111011101101000",
    "1111100010111011",
    "1111101000110010",
    "1111101111001010",
    "1111110101111111",
    "1111111101001110",
    "1111111011001101",
    "1111110011011110",
    "1111101011110000",
    "1111100100010000",
    "1111011101001110",
    "1111010110110010",
    "1111010001001101",
    "1111001100100000",
    "1111001000110000",
    "1111000101111100",
    "1111000100000011",
    "1111000011000000",
    "1111000010101001",
    "1111000010111011",
    "1111000011101001",
    "1111000100101110",
    "1111000110000100",
    "1111000111101010",
    "1111001001100111",
    "1111001100000001",
    "1111001111001000",
    "1111010011000110",
    "1111011000000011",
    "1111011101110010",
    "1111100100000110",
    "1111101010100101",
    "1111110000110001",
    "1111110110010101",
    "1111111011000110",
    "1111111111000000",
    "1111111101110010",
    "1111111011001100",
    "1111111001000101",
    "1111110111011100",
    "1111110110010100",
    "1111110101110110",
    "1111110110000100",
    "1111110111000100",
    "1111111000101111",
    "1111111010111110",
    "1111111101100011",
    "1111111111101001",
    "1111111100110110",
    "1111111010000101",
    "1111110111010100",
    "1111110100011101",
    "1111110001010101",
    "1111101101110001",
    "1111101001100111",
    "1111100100110001",
    "1111011111001101",
    "1111011001000001",
    "1111010010010010",
    "1111001011001001",
    "1111000011101001",
    "1110111011110011",
    "1110110011110100",
    "1110101011111101",
    "1110100100101001",
    "1110011110011001",
    "1110011001101011",
    "1110010110101101",
    "1110010101011101",
    "1110010101100010",
    "1110010110011101",
    "1110010111101101",
    "1110011000111100",
    "1110011010000100",
    "1110011011001010",
    "1110011100011100",
    "1110011110000101",
    "1110100000001111",
    "1110100010111011",
    "1110100110000110",
    "1110101001101111",
    "1110101101110000",
    "1110110010000010",
    "1110110110011000",
    "1110111010100011",
    "1110111110001100",
    "1111000000111001",
    "1111000010010101",
    "1111000010010000",
    "1111000000100100",
    "1110111101011100",
    "1110111001010101",
    "1110110100110011",
    "1110110000100011",
    "1110101101001111",
    "1110101011010011",
    "1110101010111000",
    "1110101100000001",
    "1110101110011110",
    "1110110010000011",
    "1110110110100101",
    "1110111011110111",
    "1111000001110110",
    "1111001000011110",
    "1111001111101001",
    "1111010111001110",
    "1111011110111010",
    "1111100110010011",
    "1111101100111111",
    "1111110010100111",
    "1111110110111000",
    "1111111001100111",
    "1111111010111000",
    "1111111010110110",
    "1111111001110101",
    "1111111000010010",
    "1111110110101010",
    "1111110101100011",
    "1111110101011100",
    "1111110110110000",
    "1111111001101000",
    "1111111101111111",
    "1111111100011101",
    "1111110110010100",
    "1111110000001000",
    "1111101010011111",
    "1111100101101110",
    "1111100001111110",
    "1111011111001111",
    "1111011101010001",
    "1111011011110111",
    "1111011010101111",
    "1111011001110000",
    "1111011000111100",
    "1111011000010011",
    "1111010111111010",
    "1111010111111010",
    "1111011000010110",
    "1111011001001100",
    "1111011010011011",
    "1111011011111010",
    "1111011101100000",
    "1111011110111011",
    "1111011111111101",
    "1111100000011001",
    "1111011111111111",
    "1111011110101101",
    "1111011100101000",
    "1111011010000001",
    "1111010111010000",
    "1111010100110001",
    "1111010010111001",
    "1111010001111110",
    "1111010010000101",
    "1111010011001111",
    "1111010101010000",
    "1111010111111111",
    "1111011011001100",
    "1111011110101011",
    "1111100010010111",
    "1111100110001110",
    "1111101010011100",
    "1111101111001010",
    "1111110100101001",
    "1111111011001001",
    "1111111101000010",
    "1111110011111011",
    "1111101001101011",
    "1111011110110110",
    "1111010100010010",
    "1111001010111111",
    "1111000011110100",
    "1110111111010010",
    "1110111101100001",
    "1110111110000111",
    "1111000000010111",
    "1111000011100010",
    "1111000111000011",
    "1111001010100010",
    "1111001101101110",
    "1111010000100110",
    "1111010011000001",
    "1111010100111001",
    "1111010101111110",
    "1111010110000100",
    "1111010101000000",
    "1111010010110001",
    "1111001111011110",
    "1111001011011000",
    "1111000110101101",
    "1111000001111000",
    "1110111101000101",
    "1110111000101010",
    "1110110100110011",
    "1110110001101011",
    "1110101111011010",
    "1110101110000100",
    "1110101101100100",
    "1110101101110111",
    "1110101110110001",
    "1110110000000111",
    "1110110001100110",
    "1110110011000011",
    "1110110100010011",
    "1110110101010011",
    "1110110110001000",
    "1110110110110111",
    "1110110111101111",
    "1110111000111111",
    "1110111010110111",
    "1110111101100001",
    "1111000001000101",
    "1111000101100010",
    "1111001010110111",
    "1111010000111101",
    "1111010111110001",
    "1111011111001111",
    "1111100111011000",
    "1111110000001010",
    "1111111001100000",
    "1111111100110000",
    "1111110010111101",
    "1111101001011100",
    "1111100000100110",
    "1111011000101010",
    "1111010001110011",
    "1111001011111101",
    "1111000110111111",
    "1111000010101100",
    "1110111110111000",
    "1110111011011110",
    "1110111000011101",
    "1110110101111110",
    "1110110100000001",
    "1110110010101001",
    "1110110001110011",
    "1110110001010111",
    "1110110001001101",
    "1110110001010010",
    "1110110001100111",
    "1110110010010010",
    "1110110011010111",
    "1110110100111110",
    "1110110111001101",
    "1110111010000010",
    "1110111101011011",
    "1111000001001000",
    "1111000101000000",
    "1111001000101111",
    "1111001100001100",
    "1111001111001101",
    "1111010001101110",
    "1111010011100111",
    "1111010100110100",
    "1111010101010011",
    "1111010101000011",
    "1111010100001101",
    "1111010010111110",
    "1111010001110001",
    "1111010000111001",
    "1111010000110000",
    "1111010001011110",
    "1111010011001011",
    "1111010101110100",
    "1111011001010001",
    "1111011101011001",
    "1111100010000011",
    "1111100111001011",
    "1111101100101000",
    "1111110010010010",
    "1111110111111101",
    "1111111101011010",
    "1111111101100101",
    "1111111001010010",
    "1111110101110001",
    "1111110011001001",
    "1111110001010111",
    "1111110000011011",
    "1111110000010011",
    "1111110000111101",
    "1111110010011010",
    "1111110100101100",
    "1111110111110111",
    "1111111100000000",
    "1111111110110111",
    "1111111000110010",
    "1111110001110011",
    "1111101001111100",
    "1111100001010100",
    "1111010111111110",
    "1111001110000101",
    "1111000100000000",
    "1110111010001110",
    "1110110001011001",
    "1110101010000110",
    "1110100100110001",
    "1110100001100111",
    "1110100000011110",
    "1110100000111011",
    "1110100010011111",
    "1110100100101110",
    "1110100111011000",
    "1110101010011001",
    "1110101101111111",
    "1110110010001101",
    "1110110111010000",
    "1110111101000100",
    "1111000011100010",
    "1111001010011011",
    "1111010001100001",
    "1111011000100010",
    "1111011111001111",
    "1111100101011010",
    "1111101010110010",
    "1111101111001010",
    "1111110010010110",
    "1111110100010110",
    "1111110101001100",
    "1111110100111101",
    "1111110011101110",
    "1111110001100011",
    "1111101110100000",
    "1111101010100110",
    "1111100101110110",
    "1111100000010101",
    "1111011010010001",
    "1111010011111000",
    "1111001101100001",
    "1111000111100101",
    "1111000010011101",
    "1110111110011111",
    "1110111011111000",
    "1110111010110000",
    "1110111011000100",
    "1110111100110000",
    "1110111111101100",
    "1111000011110001",
    "1111001000111010",
    "1111001110111011",
    "1111010101101010",
    "1111011100110111",
    "1111100100001010",
    "1111101011010100",
    "1111110010000110",
    "1111111000011001",
    "1111111110010001",
    "1111111100001010",
    "1111110110111001",
    "1111110001111011",
    "1111101101011011",
    "1111101001101101",
    "1111100111000111",
    "1111100110000000",
    "1111100110100001",
    "1111101000110101",
    "1111101100110101",
    "1111110010011001",
    "1111111001010100",
    "1111111110101111",
    "1111110110010010",
    "1111101101110011",
    "1111100101110100",
    "1111011110110110",
    "1111011001001011",
    "1111010100110110",
    "1111010001101011",
    "1111001111010010",
    "1111001101010110",
    "1111001011101101",
    "1111001010010001",
    "1111001001001011",
    "1111001000100101",
    "1111001000101100",
    "1111001001100010",
    "1111001011000110",
    "1111001101010100",
    "1111010000000010",
    "1111010011000000",
    "1111010110000011",
    "1111011000111111",
    "1111011011110000",
    "1111011110001101",
    "1111100000011100",
    "1111100010100100",
    "1111100100101111",
    "1111100111001110",
    "1111101010010000",
    "1111101110000001",
    "1111110010100110",
    "1111110111111111",
    "1111111110000000",
    "1111111011100101",
    "1111110101010001",
    "1111101111100101",
    "1111101011000110",
    "1111101000011001",
    "1111100111111100",
    "1111101001111100",
    "1111101110011010",
    "1111110100111101",
    "1111111100111111",
    "1111111010001101",
    "1111110001011111",
    "1111101001100000",
    "1111100010110011",
    "1111011101100110",
    "1111011010000110",
    "1111011000010000",
    "1111010111111111",
    "1111011001001100",
    "1111011011110000",
    "1111011111100011",
    "1111100100011100",
    "1111101010010001",
    "1111110000111000",
    "1111110111111011",
    "1111111111000011",
    "1111111010000110",
    "1111110100000000",
    "1111101110111111",
    "1111101011010110",
    "1111101001001010",
    "1111101000011010",
    "1111101000111001",
    "1111101010010110",
    "1111101100011000",
    "1111101110100101",
    "1111110000100100",
    "1111110001111110",
    "1111110010100110",
    "1111110010010111",
    "1111110001010010",
    "1111101111100010",
    "1111101101010100",
    "1111101010110100",
    "1111101000001100",
    "1111100101100010",
    "1111100010111001",
    "1111100000001101",
    "1111011101010100",
    "1111011010000110",
    "1111010110010010",
    "1111010001101110",
    "1111001100010100",
    "1111000110000011",
    "1110111111000000",
    "1110110111011011",
    "1110101111101000",
    "1110100111111001",
    "1110100000100011",
    "1110011001101111",
    "1110010011100100",
    "1110001101111111",
    "1110001000111010",
    "1110000100010000",
    "1101111111111011",
    "1101111011111010",
    "1101111000010001",
    "1101110101000101",
    "1101110010011101",
    "1101110000100100",
    "1101101111100001",
    "1101101111011111",
    "1101110000100111",
    "1101110011000011",
    "1101110110110110",
    "1101111100000101",
    "1110000010110001",
    "1110001010110000",
    "1110010011111000",
    "1110011101110010",
    "1110101000001011",
    "1110110010101001",
    "1110111100110101",
    "1111000110011010",
    "1111001111000111",
    "1111010110110111",
    "1111011101101001",
    "1111100011100001",
    "1111101000100011",
    "1111101100110111",
    "1111110000100100",
    "1111110011101111",
    "1111110110011110",
    "1111111000111010",
    "1111111011001001",
    "1111111101001011",
    "1111111111000101",
    "1111111111001011",
    "1111111101101100",
    "1111111100011010",
    "1111111011010111",
    "1111111010100010",
    "1111111001111000",
    "1111111001011000",
    "1111111001000101",
    "1111111000111111",
    "1111111001000101",
    "1111111001010111",
    "1111111001110001",
    "1111111010001101",
    "1111111010100100",
    "1111111010110100",
    "1111111010111001",
    "1111111010110110",
    "1111111010101100",
    "1111111010011011",
    "1111111010000111",
    "1111111001110001",
    "1111111001010111",
    "1111111000111010",
    "1111111000011001",
    "1111110111110011",
    "1111110111001010",
    "1111110110100011",
    "1111110110000111",
    "1111110101111101",
    "1111110110010000",
    "1111110111000110",
    "1111111000100001",
    "1111111010011110",
    "1111111100111001",
    "1111111111100111",
    "1111111101011011",
    "1111111010100000",
    "1111110111101101",
    "1111110101001011",
    "1111110011000101",
    "1111110001100010",
    "1111110000101000",
    "1111110000011011",
    "1111110000111100",
    "1111110010000110",
    "1111110011110010",
    "1111110101110111",
    "1111111000001000",
    "1111111010010101",
    "1111111100001111",
    "1111111101101001",
    "1111111110010100",
    "1111111110001011",
    "1111111101001010",
    "1111111011010101",
    "1111111000110011",
    "1111110101110001",
    "1111110010011111",
    "1111101111001101",
    "1111101100001101",
    "1111101001101000",
    "1111100111100011",
    "1111100101111001",
    "1111100100011000",
    "1111100010101110",
    "1111100000100100",
    "1111011101101011",
    "1111011001111101",
    "1111010101011111",
    "1111010000011010",
    "1111001010111101",
    "1111000101011000",
    "1110111111110101",
    "1110111010011110",
    "1110110101011011",
    "1110110000110110",
    "1110101100110010",
    "1110101001010110",
    "1110100110100101",
    "1110100100100010",
    "1110100011001011",
    "1110100010100001",
    "1110100010011111",
    "1110100011000101",
    "1110100100010010",
    "1110100110000001",
    "1110101000010011",
    "1110101011000001",
    "1110101110001010",
    "1110110001101011",
    "1110110101100101",
    "1110111001111010",
    "1110111110110000",
    "1111000100000101",
    "1111001001110101",
    "1111001111111101",
    "1111010110001110",
    "1111011100011110",
    "1111100010011001",
    "1111100111101110",
    "1111101100010111",
    "1111110000001110",
    "1111110011010011",
    "1111110101101101",
    "1111110111100000",
    "1111111000110000",
    "1111111001011111",
    "1111111001101110",
    "1111111001011111",
    "1111111000111100",
    "1111111000010101",
    "1111110111111111",
    "1111111000010000",
    "1111111001011100",
    "1111111011110010",
    "1111111111011010",
    "1111111011101010",
    "1111110101100101",
    "1111101110100101",
    "1111100110111011",
    "1111011111000010",
    "1111010111010110",
    "1111010000011010",
    "1111001010100110",
    "1111000110010011",
    "1111000011100110",
    "1111000010011100",
    "1111000010100010",
    "1111000011100100",
    "1111000101000110",
    "1111000110110110",
    "1111001000100000",
    "1111001001111100",
    "1111001010111111",
    "1111001011100000",
    "1111001011011000",
    "1111001010011001",
    "1111001000100000",
    "1111000101101001",
    "1111000001110110",
    "1110111101010100",
    "1110111000010011",
    "1110110011001101",
    "1110101110011001",
    "1110101010010011",
    "1110100111010101",
    "1110100101110100",
    "1110100101111100",
    "1110100111110100",
    "1110101011010011",
    "1110110000001010",
    "1110110110000000",
    "1110111100010001",
    "1111000010010111",
    "1111000111101101",
    "1111001011111100",
    "1111001110110011",
    "1111010000010100",
    "1111010000101110",
    "1111010000010101",
    "1111001111011111",
    "1111001110011011",
    "1111001101010010",
    "1111001100001010",
    "1111001011000010",
    "1111001001111001",
    "1111001000101000",
    "1111000111001011",
    "1111000101011111",
    "1111000011011101",
    "1111000001001101",
    "1110111110110110",
    "1110111100101101",
    "1110111011000110",
    "1110111010010011",
    "1110111010011110",
    "1110111011100000",
    "1110111101001001",
    "1110111111000010",
    "1111000000110011",
    "1111000010001000",
    "1111000010110011",
    "1111000010101110",
    "1111000001111110",
    "1111000000101001",
    "1110111110111000",
    "1110111100110101",
    "1110111010101011",
    "1110111000101111",
    "1110110111010001",
    "1110110110100101",
    "1110110111000001",
    "1110111000101100",
    "1110111011101000",
    "1110111111101001",
    "1111000100010011",
    "1111001001001011",
    "1111001101101011",
    "1111010001011010",
    "1111010100001000",
    "1111010101110001",
    "1111010110011000",
    "1111010110001000",
    "1111010101001101",
    "1111010011110001",
    "1111010001111001",
    "1111001111101100",
    "1111001101010100",
    "1111001010111010",
    "1111001000101101",
    "1111000110111110",
    "1111000101110111",
    "1111000101100010",
    "1111000110000000",
    "1111000111001101",
    "1111001001000100",
    "1111001011100000",
    "1111001110010111",
    "1111010001100110",
    "1111010101000011",
    "1111011000100000",
    "1111011011110111",
    "1111011110111011",
    "1111100001110001",
    "1111100100011100",
    "1111100111000110",
    "1111101001111100",
    "1111101101000011",
    "1111110000011100",
    "1111110100000100",
    "1111110111110011",
    "1111111011011110",
    "1111111110111011",
    "1111111101111011",
    "1111111011010110",
    "1111111001011011",
    "1111111000010001",
    "1111110111111111",
    "1111111000100100",
    "1111111001111101",
    "1111111100000100",
    "1111111110110001",
    "1111111110000001",
    "1111111010011100",
    "1111110110100001",
    "1111110010010101",
    "1111101101111100",
    "1111101001011111",
    "1111100101000101",
    "1111100000110110",
    "1111011100111010",
    "1111011001011000",
    "1111010110010101",
    "1111010011110110",
    "1111010001111101",
    "1111010000100110",
    "1111001111110011",
    "1111001111011010",
    "1111001111010111",
    "1111001111101000",
    "1111010000000111",
    "1111010000111000",
    "1111010001111011",
    "1111010011010011",
    "1111010101000110",
    "1111010111010110",
    "1111011010000111",
    "1111011101011001",
    "1111100001001100",
    "1111100101010111",
    "1111101001110100",
    "1111101110011110",
    "1111110011001110",
    "1111111000000101",
    "1111111101000110",
    "1111111101100110",
    "1111110111111101",
    "1111110001111010",
    "1111101011011101",
    "1111100100101100",
    "1111011101110000",
    "1111010110111011",
    "1111010000011100",
    "1111001010101011",
    "1111000101110110",
    "1111000010000101",
    "1110111111011010",
    "1110111101110010",
    "1110111100111111",
    "1110111100110111",
    "1110111101010100",
    "1110111110010001",
    "1110111111101100",
    "1111000001101100",
    "1111000100010101",
    "1111000111100101",
    "1111001011011110",
    "1111001111111010",
    "1111010100110011",
    "1111011010000001",
    "1111011111011110",
    "1111100100111100",
    "1111101010010110",
    "1111101111011100",
    "1111110100000011",
    "1111110111111110",
    "1111111011000011",
    "1111111101010011",
    "1111111110110000",
    "1111111111100011",
    "1111111111111000",
    "1111111111111000",
    "1111111111101000",
    "1111111111001001",
    "1111111110011001",
    "1111111101010010",
    "1111111011110100",
    "1111111001111110",
    "1111110111110100",
    "1111110101010111",
    "1111110010101001",
    "1111101111101000",
    "1111101100010000",
    "1111101000011110",
    "1111100100001110",
    "1111011111011110",
    "1111011010001110",
    "1111010100011111",
    "1111001110010001",
    "1111000111100111",
    "1111000000100011",
    "1110111001000111",
    "1110110001100001",
    "1110101001111100",
    "1110100010110011",
    "1110011100011100",
    "1110010111010101",
    "1110010011101100",
    "1110010001101100",
    "1110010001001111",
    "1110010010000101",
    "1110010011111011",
    "1110010110010110",
    "1110011001000110",
    "1110011011111100",
    "1110011110110110",
    "1110100001111001",
    "1110100101001101",
    "1110101000110100",
    "1110101100101110",
    "1110110000110101",
    "1110110100110011",
    "1110111000001110",
    "1110111010110000",
    "1110111100000010",
    "1110111011110111",
    "1110111010010011",
    "1110110111100111",
    "1110110100010010",
    "1110110000111011",
    "1110101110001100",
    "1110101100100101",
    "1110101100011100",
    "1110101101111111",
    "1110110001001000",
    "1110110101101001",
    "1110111011001111",
    "1111000001100110",
    "1111001000010000",
    "1111001110111010",
    "1111010101001000",
    "1111011010100101",
    "1111011111000101",
    "1111100010011111",
    "1111100100110111",
    "1111100110011111",
    "1111100111101011",
    "1111101000110110",
    "1111101010010010",
    "1111101100001101",
    "1111101110101010",
    "1111110001100111",
    "1111110100111010",
    "1111111000011001",
    "1111111011111011",
    "1111111111011111",
    "1111111100110111",
    "1111111001000111",
    "1111110101000111",
    "1111110000110011",
    "1111101100010000",
    "1111100111101011",
    "1111100011010011",
    "1111011111011110",
    "1111011100010100",
    "1111011010000010",
    "1111011000100011",
    "1111010111110001",
    "1111010111100010",
    "1111010111101010",
    "1111010111111111",
    "1111011000011011",
    "1111011000110101",
    "1111011001001011",
    "1111011001011000",
    "1111011001011000",
    "1111011001001001",
    "1111011000101100",
    "1111011000000001",
    "1111010111001000",
    "1111010110000001",
    "1111010100101110",
    "1111010011001111",
    "1111010001100110",
    "1111001111111010",
    "1111001110001100",
    "1111001100100110",
    "1111001011010011",
    "1111001010011000",
    "1111001010000010",
    "1111001010011011",
    "1111001011100110",
    "1111001101101101",
    "1111010000101110",
    "1111010100101100",
    "1111011001100010",
    "1111011111001000",
    "1111100101010010",
    "1111101011110000",
    "1111110010011000",
    "1111111001000001",
    "1111111111101011",
    "1111111001100010",
    "1111110010101101",
    "1111101011111000",
    "1111100101010010",
    "1111011111010001",
    "1111011010001100",
    "1111010110011011",
    "1111010100000011",
    "1111010010111101",
    "1111010010111000",
    "1111010011100010",
    "1111010100101010",
    "1111010110000001",
    "1111010111100000",
    "1111011001000100",
    "1111011010100011",
    "1111011011110011",
    "1111011100100011",
    "1111011100100000",
    "1111011011011001",
    "1111011001001011",
    "1111010101111001",
    "1111010001110011",
    "1111001101001111",
    "1111001000100010",
    "1111000100000000",
    "1110111111110110",
    "1110111100001010",
    "1110111000111111",
    "1110110110010010",
    "1110110100000000",
    "1110110010000010",
    "1110110000001111",
    "1110101110100100",
    "1110101100111101",
    "1110101011011001",
    "1110101001111100",
    "1110101000101101",
    "1110100111110101",
    "1110100111011011",
    "1110100111100010",
    "1110101000001110",
    "1110101001011110",
    "1110101011010110",
    "1110101101110011",
    "1110110000111101",
    "1110110100110100",
    "1110111001011001",
    "1110111110101110",
    "1111000100101111",
    "1111001011010100",
    "1111010010011010",
    "1111011001110111",
    "1111100001100111",
    "1111101001101100",
    "1111110010000100",
    "1111111010101101",
    "1111111100011010",
    "1111110011100100",
    "1111101010111001",
    "1111100010101110",
    "1111011011001010",
    "1111010100011100",
    "1111001110011111",
    "1111001001010110",
    "1111000100111011",
    "1111000001001000",
    "1110111101111101",
    "1110111011010100",
    "1110111001001001",
    "1110110111011011",
    "1110110110000110",
    "1110110101001000",
    "1110110100100101",
    "1110110100100010",
    "1110110101000011",
    "1110110110001110",
    "1110111000000110",
    "1110111010101111",
    "1110111110000101",
    "1111000010001010",
    "1111000110110001",
    "1111001011101010",
    "1111010000100011",
    "1111010101000110",
    "1111011000111010",
    "1111011011101011",
    "1111011101000111",
    "1111011101001111",
    "1111011100001110",
    "1111011010011011",
    "1111011000011010",
    "1111010110100101",
    "1111010101011011",
    "1111010101001000",
    "1111010101101100",
    "1111010111000110",
    "1111011001010011",
    "1111011100010001",
    "1111100000000011",
    "1111100100101100",
    "1111101010001100",
    "1111110000011000",
    "1111110110111101",
    "1111111101100101",
    "1111111100001010",
    "1111110110101011",
    "1111110010001011",
    "1111101110101111",
    "1111101100010111",
    "1111101010111100",
    "1111101010011001",
    "1111101010101000",
    "1111101011100110",
    "1111101101010010",
    "1111101111101101",
    "1111110010111101",
    "1111110111000111",
    "1111111100010001",
    "1111111101100000",
    "1111110110010100",
    "1111101110001011",
    "1111100101001110",
    "1111011011100101",
    "1111010001011111",
    "1111000111010101",
    "1110111101101000",
    "1110110101000011",
    "1110101110001111",
    "1110101001101000",
    "1110100111011010",
    "1110100111010101",
    "1110101000111111",
    "1110101011111000",
    "1110101111100001",
    "1110110011100110",
    "1110110111111110",
    "1110111100100011",
    "1111000001011001",
    "1111000110011010",
    "1111001011011101",
    "1111010000011100",
    "1111010101001011",
    "1111011001100101",
    "1111011101100110",
    "1111100001001010",
    "1111100100001101",
    "1111100110101100",
    "1111101000100100",
    "1111101001110011",
    "1111101010011011",
    "1111101010011101",
    "1111101001111000",
    "1111101000101000",
    "1111100110101000",
    "1111100011101111",
    "1111011111111101",
    "1111011011010011",
    "1111010101111001",
    "1111010000000011",
    "1111001010001001",
    "1111000100100000",
    "1110111111011100",
    "1110111011001001",
    "1110110111101101",
    "1110110101001000",
    "1110110011011101",
    "1110110010110001",
    "1110110011000110",
    "1110110100101001",
    "1110110111011011",
    "1110111011100011",
    "1111000000111011",
    "1111000111011010",
    "1111001110101001",
    "1111010110010010",
    "1111011101110101",
    "1111100100111011",
    "1111101011010101",
    "1111110000111101",
    "1111110101110111",
    "1111111010001011",
    "1111111110000010",
    "1111111110011101",
    "1111111011011011",
    "1111111000111010",
    "1111110111000110",
    "1111110110001000",
    "1111110110000011",
    "1111110110111100",
    "1111111000110010",
    "1111111011100111",
    "1111111111011110",
    "1111111011100011",
    "1111110101100010",
    "1111101110100010",
    "1111100110111010",
    "1111011111000111",
    "1111010111101101",
    "1111010001001111",
    "1111001100000101",
    "1111001000010101",
    "1111000101110100",
    "1111000100001110",
    "1111000011001011",
    "1111000010010101",
    "1111000001101011",
    "1111000001001100",
    "1111000001000111",
    "1111000001101001",
    "1111000010111001",
    "1111000100111011",
    "1111000111100111",
    "1111001010110101",
    "1111001110011100",
    "1111010010010111",
    "1111010110100000",
    "1111011010110100",
    "1111011111010010",
    "1111100011111001",
    "1111101000100101",
    "1111101101010100",
    "1111110010000110",
    "1111110110111001",
    "1111111011101101",
    "1111111111011111",
    "1111111010111010",
    "1111110110110010",
    "1111110011011111",
    "1111110001011011",
    "1111110000111111",
    "1111110010011101",
    "1111110101111101",
    "1111111011010011",
    "1111111101110101",
    "1111110110000111",
    "1111101110001101",
    "1111100110111001",
    "1111100000110001",
    "1111011100010100",
    "1111011001101111",
    "1111011000111111",
    "1111011001110010",
    "1111011011110101",
    "1111011110110011",
    "1111100010011100",
    "1111100110100101",
    "1111101011001000",
    "1111101111111111",
    "1111110100111111",
    "1111111001111101",
    "1111111110101010",
    "1111111101000100",
    "1111111001011111",
    "1111110110101000",
    "1111110100100100",
    "1111110011010001",
    "1111110010101010",
    "1111110010100111",
    "1111110010111111",
    "1111110011100000",
    "1111110011111101",
    "1111110100000110",
    "1111110011110001",
    "1111110010111001",
    "1111110001011111",
    "1111101111101010",
    "1111101101100011",
    "1111101011010010",
    "1111101001000000",
    "1111100110110001",
    "1111100100100101",
    "1111100010011100",
    "1111100000010001",
    "1111011101111000",
    "1111011011001010",
    "1111010111111110",
    "1111010100001000",
    "1111001111100100",
    "1111001010001100",
    "1111000100000011",
    "1110111101001100",
    "1110110101110010",
    "1110101110000111",
    "1110100110011101",
    "1110011111001100",
    "1110011000100101",
    "1110010010110110",
    "1110001110000010",
    "1110001010000001",
    "1110000110101000",
    "1110000011100111",
    "1110000000110001",
    "1101111110001001",
    "1101111011110010",
    "1101111001111010",
    "1101111000110010",
    "1101111000100101",
    "1101111001011001",
    "1101111011001110",
    "1101111101111010",
    "1110000001010111",
    "1110000101011010",
    "1110001010000001",
    "1110001111000101",
    "1110010100100111",
    "1110011010100010",
    "1110100000101110",
    "1110100110111111",
    "1110101101001010",
    "1110110010111110",
    "1110111000010110",
    "1110111101001111",
    "1111000001110100",
    "1111000110010000",
    "1111001010110000",
    "1111001111011110",
    "1111010100011000",
    "1111011001011001",
    "1111011110010100",
    "1111100010110110",
    "1111100110110011",
    "1111101010000110",
    "1111101100110000",
    "1111101110111000",
    "1111110000101100",
    "1111110010010100",
    "1111110011111001",
    "1111110101011011",
    "1111110110111000",
    "1111111000001011",
    "1111111001001111",
    "1111111010000011",
    "1111111010100101",
    "1111111010111000",
    "1111111011000010",
    "1111111011001000",
    "1111111011010001",
    "1111111011100111",
    "1111111100010101",
    "1111111101100000",
    "1111111111010001",
    "1111111110010110",
    "1111111011100000",
    "1111111000010011",
    "1111110101000010",
    "1111110001111111",
    "1111101111100000",
    "1111101101110111",
    "1111101101010001",
    "1111101101110011",
    "1111101111011000",
    "1111110001110100",
    "1111110100110110",
    "1111111000001100",
    "1111111011100110",
    "1111111110111001",
    "1111111101111101",
    "1111111011000010",
    "1111111000010001",
    "1111110101101000",
    "1111110011001010",
    "1111110000111100",
    "1111101111000111",
    "1111101101110011",
    "1111101101000111",
    "1111101101000110",
    "1111101101101110",
    "1111101110110111",
    "1111110000011000",
    "1111110010000011",
    "1111110011110001",
    "1111110101011011",
    "1111110110111111",
    "1111111000011110",
    "1111111001111001",
    "1111111011010001",
    "1111111100100110",
    "1111111101110101",
    "1111111110111110",
    "1111111111111101",
    "1111111111001100",
    "1111111110100111",
    "1111111110010101",
    "1111111110100001",
    "1111111111010101",
    "1111111111000000",
    "1111111100010111",
    "1111111000101100",
    "1111110011111111",
    "1111101110011010",
    "1111101000001010",
    "1111100001100001",
    "1111011010101111",
    "1111010100000011",
    "1111001101110000",
    "1111000111111110",
    "1111000010111000",
    "1110111110011011",
    "1110111010100011",
    "1110110111001001",
    "1110110100000101",
    "1110110001010000",
    "1110101110110011",
    "1110101100110011",
    "1110101011011011",
    "1110101010110010",
    "1110101010111100",
    "1110101011110011",
    "1110101101010100",
    "1110101111010010",
    "1110110001101011",
    "1110110100011000",
    "1110110111100000",
    "1110111011000110",
    "1110111111001101",
    "1111000011111001",
    "1111001001000110",
    "1111001110101001",
    "1111010100011000",
    "1111011010000001",
    "1111011111010111",
    "1111100100001110",
    "1111101000100001",
    "1111101100001100",
    "1111101111010001",
    "1111110001110101",
    "1111110011111110",
    "1111110101110000",
    "1111110111010010",
    "1111111000100111",
    "1111111001110000",
    "1111111010101110",
    "1111111011100010",
    "1111111100001100",
    "1111111100110001",
    "1111111101011010",
    "1111111110010101",
    "1111111111110100",
    "1111111101110100",
    "1111111010011110",
    "1111110110000000",
    "1111110000100001",
    "1111101010010001",
    "1111100011101010",
    "1111011101001100",
    "1111010111011011",
    "1111010010111000",
    "1111001111111000",
    "1111001110101101",
    "1111001111001111",
    "1111010001001100",
    "1111010011111100",
    "1111010110110111",
    "1111011001001100",
    "1111011010010110",
    "1111011010000001",
    "1111011000000001",
    "1111010100011101",
    "1111001111100011",
    "1111001001100000",
    "1111000010100111",
    "1110111011001001",
    "1110110011011101",
    "1110101100000001",
    "1110100101011000",
    "1110100000000111",
    "1110011100101110",
    "1110011011100001",
    "1110011100101000",
    "1110011111110011",
    "1110100100101110",
    "1110101010110111",
    "1110110001110011",
    "1110111001000010",
    "1111000000001100",
    "1111000110110010",
    "1111001100011110",
    "1111010000111011",
    "1111010011111110",
    "1111010101100100",
    "1111010101110111",
    "1111010101001011",
    "1111010011110100",
    "1111010010001010",
    "1111010000011110",
    "1111001110110110",
    "1111001101011100",
    "1111001100010001",
    "1111001011011000",
    "1111001010101011",
    "1111001010001100",
    "1111001001110101",
    "1111001001011101",
    "1111001000111100",
    "1111001000010000",
    "1111000111010110",
    "1111000110010101",
    "1111000101010000",
    "1111000100010010",
    "1111000011100001",
    "1111000011000000",
    "1111000010110001",
    "1111000010101110",
    "1111000010110100",
    "1111000010111101",
    "1111000011000000",
    "1111000011000000",
    "1111000010111011",
    "1111000010110110",
    "1111000010111000",
    "1111000011000011",
    "1111000011011010",
    "1111000011111001",
    "1111000100011101",
    "1111000101000000",
    "1111000101100000",
    "1111000110000001",
    "1111000110101000",
    "1111000111100000",
    "1111001000101010",
    "1111001010000100",
    "1111001011100001",
    "1111001100110111",
    "1111001101110000",
    "1111001110000111",
    "1111001101110011",
    "1111001100111000",
    "1111001011011101",
    "1111001001101101",
    "1111000111110101",
    "1111000110000110",
    "1111000100101110",
    "1111000011110110",
    "1111000011101100",
    "1111000100011000",
    "1111000101111100",
    "1111001000100000",
    "1111001100000010",
    "1111010000100100",
    "1111010101110110",
    "1111011011101000",
    "1111100001100010",
    "1111100111001000",
    "1111101100000011",
    "1111110000000110",
    "1111110011010000",
    "1111110101101000",
    "1111110111100001",
    "1111111001001001",
    "1111111010110000",
    "1111111100100000",
    "1111111110011111",
    "1111111111010011",
    "1111111100111110",
    "1111111010100100",
    "1111111000001010",
    "1111110101110110",
    "1111110011101101",
    "1111110001110010",
    "1111110000001010",
    "1111101110111111",
    "1111101110011000",
    "1111101110100100",
    "1111101111110011",
    "1111110010011000",
    "1111110110100010",
    "1111111100011101",
    "1111111011111001",
    "1111110010111000",
    "1111101001001000",
    "1111011111011100",
    "1111010110101100",
    "1111001111011111",
    "1111001010010011",
    "1111000111000110",
    "1111000101100100",
    "1111000101001110",
    "1111000101101001",
    "1111000110011000",
    "1111000111010011",
    "1111001000011010",
    "1111001001101111",
    "1111001011011001",
    "1111001101011110",
    "1111001111111010",
    "1111010010100111",
    "1111010101100010",
    "1111011000100011",
    "1111011011101010",
    "1111011110101110",
    "1111100001110000",
    "1111100100101110",
    "1111100111101001",
    "1111101010100100",
    "1111101101100101",
    "1111110000111000",
    "1111110100100011",
    "1111111000110011",
    "1111111101101001",
    "1111111100111001",
    "1111110111000100",
    "1111110001000101",
    "1111101011010100",
    "1111100110000110",
    "1111100001101100",
    "1111011110001111",
    "1111011011101011",
    "1111011001110111",
    "1111011000100010",
    "1111010111011000",
    "1111010110001110",
    "1111010100111110",
    "1111010011100110",
    "1111010010001011",
    "1111010000111000",
    "1111001111110101",
    "1111001111000101",
    "1111001110110101",
    "1111001111001111",
    "1111010000100001",
    "1111010010111011",
    "1111010110101101",
    "1111011011111111",
    "1111100010101100",
    "1111101010011111",
    "1111110010110011",
    "1111111010111101",
    "1111111101110000",
    "1111110111111100",
    "1111110011110100",
    "1111110001011000",
    "1111110000010110",
    "1111110000010110",
    "1111110001000001",
    "1111110010000101",
    "1111110011011010",
    "1111110100111101",
    "1111110110101111",
    "1111111000110000",
    "1111111011000000",
    "1111111101011001",
    "1111111111111001",
    "1111111101100011",
    "1111111011000000",
    "1111111000011010",
    "1111110101101011",
    "1111110010101001",
    "1111101111001011",
    "1111101011000111",
    "1111100110010101",
    "1111100000110001",
    "1111011010011101",
    "1111010011011111",
    "1111001100000010",
    "1111000100010101",
    "1110111100100101",
    "1110110100111110",
    "1110101101110011",
    "1110100111010110",
    "1110100001111001",
    "1110011101101110",
    "1110011011000110",
    "1110011010000100",
    "1110011010101011",
    "1110011100101101",
    "1110011111111011",
    "1110100011111001",
    "1110101000001110",
    "1110101100010111",
    "1110101111111101",
    "1110110010100010",
    "1110110011111001",
    "1110110011111110",
    "1110110010111001",
    "1110110000111011",
    "1110101110011111",
    "1110101100000001",
    "1110101001110101",
    "1110101000001011",
    "1110100111000110",
    "1110100110100111",
    "1110100110100101",
    "1110100110111110",
    "1110100111101010",
    "1110101000110010",
    "1110101010011110",
    "1110101100111100",
    "1110110000010111",
    "1110110100111001",
    "1110111010011110",
    "1111000000110110",
    "1111000111101100",
    "1111001110011011",
    "1111010100100100",
    "1111011001101010",
    "1111011101011110",
    "1111100000000000",
    "1111100001011010",
    "1111100010000010",
    "1111100010010000",
    "1111100010011101",
    "1111100011000101",
    "1111100100010101",
    "1111100110011110",
    "1111101001100010",
    "1111101101100010",
    "1111110010001111",
    "1111110111010111",
    "1111111100100100",
    "1111111110011100",
    "1111111001111111",
    "1111110110001001",
    "1111110010111001",
    "1111110000001010",
    "1111101101110101",
    "1111101011110011",
    "1111101010000110",
    "1111101000110000",
    "1111100111110101",
    "1111100111010111",
    "1111100111010001",
    "1111100111011111",
    "1111100111111000",
    "1111101000011000",
    "1111101000111000",
    "1111101001010101",
    "1111101001101011",
    "1111101001110011",
    "1111101001100011",
    "1111101000101111",
    "1111100111001110",
    "1111100100111001",
    "1111100001110110",
    "1111011110010010",
    "1111011010100011",
    "1111010110111110",
    "1111010011111001",
    "1111010001100111",
    "1111010000001111",
    "1111001111101110",
    "1111001111111101",
    "1111010000110001",
    "1111010001111011",
    "1111010011010010",
    "1111010100110110",
    "1111010110101100",
    "1111011001000001",
    "1111011100000010",
    "1111011111111111",
    "1111100100110111",
    "1111101010101001",
    "1111110001000001",
    "1111110111100111",
    "1111111110000100",
    "1111111011111001",
    "1111110110011100",
    "1111110001011111",
    "1111101100111001",
    "1111101000100011",
    "1111100100011000",
    "1111100000011110",
    "1111011100111101",
    "1111011001111101",
    "1111010111100101",
    "1111010101110010",
    "1111010100011100",
    "1111010011011100",
    "1111010010100111",
    "1111010001111110",
    "1111010001011100",
    "1111010001000011",
    "1111010000101110",
    "1111010000011010",
    "1111001111111111",
    "1111001111010010",
    "1111001110000111",
    "1111001100010111",
    "1111001001111010",
    "1111000110101111",
    "1111000010111001",
    "1110111110100011",
    "1110111001111010",
    "1110110101010101",
    "1110110001000000",
    "1110101101001100",
    "1110101010000010",
    "1110100111100010",
    "1110100101101001",
    "1110100100001101",
    "1110100011001011",
    "1110100010011111",
    "1110100010001101",
    "1110100010011001",
    "1110100011001101",
    "1110100100110100",
    "1110100111010000",
    "1110101010100011",
    "1110101110100011",
    "1110110011000000",
    "1110110111101111",
    "1110111100011011",
    "1111000000110101",
    "1111000100110110",
    "1111001000011010",
    "1111001011100101",
    "1111001110100100",
    "1111010001100111",
    "1111010101000000",
    "1111011000111100",
    "1111011101101011",
    "1111100011010011",
    "1111101001111100",
    "1111110001100100",
    "1111111010000101",
    "1111111100101010",
    "1111110011000100",
    "1111101001100001",
    "1111100000100011",
    "1111011000100111",
    "1111010010000011",
    "1111001100111111",
    "1111001001011000",
    "1111000110111001",
    "1111000101001011",
    "1111000011110110",
    "1111000010100100",
    "1111000001001010",
    "1110111111100100",
    "1110111101110111",
    "1110111100001001",
    "1110111010100101",
    "1110111001010011",
    "1110111000011101",
    "1110111000001001",
    "1110111000011101",
    "1110111001011101",
    "1110111011000110",
    "1110111101001110",
    "1110111111101000",
    "1111000010000000",
    "1111000100001000",
    "1111000101110100",
    "1111000110111110",
    "1111000111100111",
    "1111000111111010",
    "1111001000000011",
    "1111001000010000",
    "1111001000101101",
    "1111001001100010",
    "1111001010110010",
    "1111001100100000",
    "1111001110101001",
    "1111010001010100",
    "1111010100011101",
    "1111011000010001",
    "1111011100110101",
    "1111100010000110",
    "1111101000000101",
    "1111101110100011",
    "1111110101010001",
    "1111111011111000",
    "1111111101111011",
    "1111111000100110",
    "1111110100010101",
    "1111110001010010",
    "1111101111100001",
    "1111101111000010",
    "1111101111110000",
    "1111110001101000",
    "1111110100100100",
    "1111111000100100",
    "1111111101100111",
    "1111111100010011",
    "1111110101001111",
    "1111101101010000",
    "1111100100100000",
    "1111011011001010",
    "1111010001100001",
    "1111000111111001",
    "1110111110110101",
    "1110110110110111",
    "1110110000100001",
    "1110101100001001",
    "1110101001110000",
    "1110101001001100",
    "1110101001111111",
    "1110101011101011",
    "1110101101111010",
    "1110110000011111",
    "1110110011100001",
    "1110110111001001",
    "1110111011100001",
    "1111000000101100",
    "1111000110011111",
    "1111001100100101",
    "1111010010100001",
    "1111010111111110",
    "1111011100100110",
    "1111100000010010",
    "1111100010111101",
    "1111100100101111",
    "1111100101101111",
    "1111100110001011",
    "1111100110001011",
    "1111100101110111",
    "1111100101010011",
    "1111100100011111",
    "1111100011010101",
    "1111100001101110",
    "1111011111100011",
    "1111011100101010",
    "1111011000111100",
    "1111010100010111",
    "1111001110111101",
    "1111001001000010",
    "1111000010111011",
    "1110111101000101",
    "1110111000000001",
    "1110110100000011",
    "1110110001010111",
    "1110101111111101",
    "1110101111101011",
    "1110110000010010",
    "1110110001101011",
    "1110110011101111",
    "1110110110100111",
    "1110111010100000",
    "1110111111100011",
    "1111000101111001",
    "1111001101011100",
    "1111010101111110",
    "1111011110111111",
    "1111101000000101",
    "1111110000110011",
    "1111111000110101",
    "1111111111111011",
    "1111111001111111",
    "1111110101000110",
    "1111110001011001",
    "1111101110111111",
    "1111101101111000",
    "1111101110000101",
    "1111101111100001",
    "1111110010000010",
    "1111110101011011",
    "1111111001011111",
    "1111111101111110",
    "1111111101010011",
    "1111111000101001",
    "1111110100001011",
    "1111101111111110",
    "1111101100000010",
    "1111101000010010",
    "1111100100100100",
    "1111100000110000",
    "1111011100101110",
    "1111011000100011",
    "1111010100010101",
    "1111010000001101",
    "1111001100011100",
    "1111001001001100",
    "1111000110101000",
    "1111000100110110",
    "1111000011110110",
    "1111000011101001",
    "1111000100001010",
    "1111000101011000",
    "1111000111010101",
    "1111001010000010",
    "1111001101100011",
    "1111010001111011",
    "1111010111001001",
    "1111011101000010",
    "1111100011011000",
    "1111101001110110",
    "1111110000000101",
    "1111110101110000",
    "1111111010101100",
    "1111111110101110",
    "1111111110001101",
    "1111111100001100",
    "1111111011001111",
    "1111111011010111",
    "1111111100100000",
    "1111111110100100",
    "1111111110101011",
    "1111111011100101",
    "1111111000011010",
    "1111110101011011",
    "1111110010110100",
    "1111110000101000",
    "1111101110111000",
    "1111101101011011",
    "1111101100001110",
    "1111101011001011",
    "1111101010010110",
    "1111101001110100",
    "1111101001110001",
    "1111101010011000",
    "1111101011110001",
    "1111101110000001",
    "1111110001000100",
    "1111110100110001",
    "1111111000110111",
    "1111111101000111",
    "1111111110101101",
    "1111111010110111",
    "1111110111011110",
    "1111110100100110",
    "1111110010010000",
    "1111110000011110",
    "1111101111010010",
    "1111101110101101",
    "1111101110101110",
    "1111101111010001",
    "1111110000010010",
    "1111110001100011",
    "1111110010111010",
    "1111110100001111",
    "1111110101011001",
    "1111110110010101",
    "1111110111000001",
    "1111110111011010",
    "1111110111011011",
    "1111110110111010",
    "1111110101101011",
    "1111110011100110",
    "1111110000100101",
    "1111101100101000",
    "1111100111110101",
    "1111100010010100",
    "1111011100001110",
    "1111010101101001",
    "1111001110101011",
    "1111000111010011",
    "1110111111100100",
    "1110110111100111",
    "1110101111100011",
    "1110100111101100",
    "1110100000010001",
    "1110011001011110",
    "1110010011011101",
    "1110001110001010",
    "1110001001011101",
    "1110000101010011",
    "1110000001101001",
    "1101111110011110",
    "1101111011111010",
    "1101111010000111",
    "1101111001010000",
    "1101111001010101",
    "1101111010011011",
    "1101111100011100",
    "1101111111010010",
    "1110000010101111",
    "1110000110101100",
    "1110001010111100",
    "1110001111011001",
    "1110010100000000",
    "1110011000101010",
    "1110011101010111",
    "1110100010000101",
    "1110100110101101",
    "1110101011001110",
    "1110101111011111",
    "1110110011100010",
    "1110110111011011",
    "1110111011010001",
    "1110111111001111",
    "1111000011100110",
    "1111001000100010",
    "1111001110001100",
    "1111010100100000",
    "1111011011011001",
    "1111100010011010",
    "1111101001000101",
    "1111101110111100",
    "1111110011100111",
    "1111110110111100",
    "1111111001000000",
    "1111111010000011",
    "1111111010011011",
    "1111111010100010",
    "1111111010100100",
    "1111111010101101",
    "1111111011000000",
    "1111111011011010",
    "1111111011111010",
    "1111111100011101",
    "1111111101000110",
    "1111111101110110",
    "1111111110110100",
    "1111111111110110",
    "1111111110000111",
    "1111111011111001",
    "1111111001000111",
    "1111110101110110",
    "1111110010001100",
    "1111101110011010",
    "1111101010110010",
    "1111100111101010",
    "1111100101010111",
    "1111100100000110",
    "1111100100000000",
    "1111100100111110",
    "1111100110111000",
    "1111101001011100",
    "1111101100011000",
    "1111101111011101",
    "1111110010011111",
    "1111110101011000",
    "1111111000000110",
    "1111111010101011",
    "1111111101001110",
    "1111111111110011",
    "1111111101011100",
    "1111111010100100",
    "1111110111100011",
    "1111110100011111",
    "1111110001100001",
    "1111101110111001",
    "1111101100110001",
    "1111101011010111",
    "1111101010110010",
    "1111101011000001",
    "1111101100000010",
    "1111101101101100",
    "1111101111110111",
    "1111110010011111",
    "1111110101011101",
    "1111111000110000",
    "1111111100010101",
    "1111111111110110",
    "1111111100000001",
    "1111111000010100",
    "1111110101000011",
    "1111110010011111",
    "1111110000111010",
    "1111110000100110",
    "1111110001101010",
    "1111110100001010",
    "1111111000000001",
    "1111111101000111",
    "1111111100110001",
    "1111110110000001",
    "1111101110111111",
    "1111101000000100",
    "1111100001100111",
    "1111011011111010",
    "1111010110111111",
    "1111010010110011",
    "1111001111000010",
    "1111001011010100",
    "1111000111010101",
    "1111000010110110",
    "1110111101110101",
    "1110111000011101",
    "1110110011000001",
    "1110101101110111",
    "1110101001010110",
    "1110100101110001",
    "1110100011010111",
    "1110100010001111",
    "1110100010011010",
    "1110100011110110",
    "1110100110011000",
    "1110101001110100",
    "1110101101111010",
    "1110110010100010",
    "1110110111100000",
    "1110111100101011",
    "1111000001111101",
    "1111000111001110",
    "1111001100010011",
    "1111010000111110",
    "1111010101000110",
    "1111011000011110",
    "1111011011000100",
    "1111011100110011",
    "1111011101110111",
    "1111011110011100",
    "1111011110110101",
    "1111011111010110",
    "1111100000010101",
    "1111100010000011",
    "1111100100101100",
    "1111101000010011",
    "1111101100110010",
    "1111110001111010",
    "1111110111011010",
    "1111111101000010",
    "1111111101011011",
    "1111111000001101",
    "1111110011011000",
    "1111101111000001",
    "1111101011001110",
    "1111101000000111",
    "1111100101101111",
    "1111100100001101",
    "1111100011011000",
    "1111100011001010",
    "1111100011010000",
    "1111100011011100",
    "1111100011100001",
    "1111100011010011",
    "1111100010110110",
    "1111100010001000",
    "1111100001001010",
    "1111011111111010",
    "1111011110010111",
    "1111011100100000",
    "1111011010001100",
    "1111010111011101",
    "1111010100010000",
    "1111010000100111",
    "1111001100100101",
    "1111001000001011",
    "1111000011100100",
    "1110111110110110",
    "1110111010010011",
    "1110110110001101",
    "1110110011000000",
    "1110110001000111",
    "1110110000111011",
    "1110110010110011",
    "1110110110110001",
    "1110111100101010",
    "1111000011111100",
    "1111001011111101",
    "1111010011101111",
    "1111011010100010",
    "1111011111101100",
    "1111100011000000",
    "1111100100100010",
    "1111100100101001",
    "1111100011110001",
    "1111100010010101",
    "1111100000100011",
    "1111011110011100",
    "1111011011111101",
    "1111011000111111",
    "1111010101011111",
    "1111010001011111",
    "1111001101001010",
    "1111001000110100",
    "1111000100101100",
    "1111000001000010",
    "1110111110000101",
    "1110111011111100",
    "1110111010101010",
    "1110111010010001",
    "1110111010100101",
    "1110111011100000",
    "1110111100110000",
    "1110111110001100",
    "1110111111101001",
    "1111000001000010",
    "1111000010010100",
    "1111000011100010",
    "1111000100110011",
    "1111000110000110",
    "1111000111100010",
    "1111001001001011",
    "1111001011000001",
    "1111001101000010",
    "1111001111001010",
    "1111010001010000",
    "1111010011010000",
    "1111010101000000",
    "1111010110010110",
    "1111010111010011",
    "1111010111101111",
    "1111010111101000",
    "1111010111000011",
    "1111010101111110",
    "1111010100011101",
    "1111010010100100",
    "1111010000010101",
    "1111001101101110",
    "1111001010101111",
    "1111000111010101",
    "1111000011100100",
    "1110111111100110",
    "1110111011101101",
    "1110111000001110",
    "1110110101100100",
    "1110110100000001",
    "1110110011110110",
    "1110110101001000",
    "1110110111110101",
    "1110111011110010",
    "1111000000101110",
    "1111000110010011",
    "1111001100000101",
    "1111010001101001",
    "1111010110100010",
    "1111011010011001",
    "1111011101001001",
    "1111011110110011",
    "1111011111101011",
    "1111100000001111",
    "1111100000111011",
    "1111100010001010",
    "1111100100001011",
    "1111100110111110",
    "1111101010011111",
    "1111101110100001",
    "1111110010111000",
    "1111110111010111",
    "1111111011110001",
    "1111111111111110",
    "1111111100001010",
    "1111111000110111",
    "1111110110001011",
    "1111110100001111",
    "1111110011000110",
    "1111110010110101",
    "1111110011100011",
    "1111110101011001",
    "1111111000100101",
    "1111111101011000",
    "1111111100000000",
    "1111110011100111",
    "1111101001101110",
    "1111011111000010",
    "1111010100100010",
    "1111001011010100",
    "1111000100010010",
    "1110111111110101",
    "1110111101111010",
    "1110111101111000",
    "1110111110111101",
    "1111000000010010",
    "1111000001010111",
    "1111000001111110",
    "1111000010010010",
    "1111000010100111",
    "1111000011010011",
    "1111000100100101",
    "1111000110100100",
    "1111001001001110",
    "1111001100011100",
    "1111010000001010",
    "1111010100001011",
    "1111011000011011",
    "1111011100101101",
    "1111100000110110",
    "1111100100110011",
    "1111101000011100",
    "1111101011111000",
    "1111101111000110",
    "1111110010001111",
    "1111110101010011",
    "1111111000010110",
    "1111111011011010",
    "1111111110011110",
    "1111111110010111",
    "1111111011001011",
    "1111110111111000",
    "1111110100011110",
    "1111110000111011",
    "1111101101010000",
    "1111101001011000",
    "1111100101010011",
    "1111100000111110",
    "1111011100011110",
    "1111010111111010",
    "1111010011100100",
    "1111001111101110",
    "1111001100110011",
    "1111001011001001",
    "1111001011000010",
    "1111001100101010",
    "1111001111111011",
    "1111010100101110",
    "1111011010101011",
    "1111100001011010",
    "1111101000011010",
    "1111101111001110",
    "1111110101011001",
    "1111111010101001",
    "1111111110110011",
    "1111111110000011",
    "1111111011111000",
    "1111111010011001",
    "1111111001011010",
    "1111111000110001",
    "1111111000011010",
    "1111111000010011",
    "1111111000011110",
    "1111111000111001",
    "1111111001100001",
    "1111111010001111",
    "1111111010111111",
    "1111111011101100",
    "1111111100010111",
    "1111111101000111",
    "1111111110000110",
    "1111111111011110",
    "1111111110011110",
    "1111111011101000",
    "1111110111110011",
    "1111110010110011",
    "1111101100100011",
    "1111100101000011",
    "1111011100011110",
    "1111010011000101",
    "1111001001011001",
    "1111000000000010",
    "1110110111100101",
    "1110110000101011",
    "1110101011100110",
    "1110101000100101",
    "1110100111011011",
    "1110100111101111",
    "1110101001000110",
    "1110101010111100",
    "1110101100111100",
    "1110101110111000",
    "1110110000101100",
    "1110110010011111",
    "1110110100010101",
    "1110110110010000",
    "1110111000001100",
    "1110111010000001",
    "1110111011011101",
    "1110111100001110",
    "1110111100000111",
    "1110111010111101",
    "1110111000101111",
    "1110110101011111",
    "1110110001011001",
    "1110101100101011",
    "1110100111110001",
    "1110100010111110",
    "1110011110101110",
    "1110011011010110",
    "1110011001000100",
    "1110010111111110",
    "1110011000000100",
    "1110011001010011",
    "1110011011100000",
    "1110011110100011",
    "1110100010010010",
    "1110100110101000",
    "1110101011011110",
    "1110110000100110",
    "1110110101110110",
    "1110111010111100",
    "1110111111100100",
    "1111000011011100",
    "1111000110010101",
    "1111001000001001",
    "1111001000111010",
    "1111001000110100",
    "1111001000001110",
    "1111000111100000",
    "1111000111000100",
    "1111000111010101",
    "1111001000100101",
    "1111001011001010",
    "1111001111001111",
    "1111010100111110",
    "1111011100010100",
    "1111100101000011",
    "1111101110101101",
    "1111111000100011",
    "1111111110001010",
    "1111110110010010",
    "1111110000010101",
    "1111101100011111",
    "1111101010100110",
    "1111101010010001",
    "1111101010111100",
    "1111101100000100",
    "1111101101010011",
    "1111101110010111",
    "1111101111001010",
    "1111101111100111",
    "1111101111101011",
    "1111101111010001",
    "1111101110010100",
    "1111101100101011",
    "1111101010010111",
    "1111100111010110",
    "1111100011101110",
    "1111011111101011",
    "1111011011010110",
    "1111010111000011",
    "1111010011000001",
    "1111001111100011",
    "1111001100110111",
    "1111001011001010",
    "1111001010100110",
    "1111001011001001",
    "1111001100101110",
    "1111001111001100",
    "1111010010010010",
    "1111010101101111",
    "1111011001010001",
    "1111011100101000",
    "1111011111100110",
    "1111100010000011",
    "1111100100000000",
    "1111100101100010",
    "1111100110111000",
    "1111101000010010",
    "1111101001111111",
    "1111101100001101",
    "1111101111000110",
    "1111110010101100",
    "1111110111000001",
    "1111111100000010",
    "1111111110010011",
    "1111111000010000",
    "1111110010000100",
    "1111101100000111",
    "1111100110111001",
    "1111100010110011",
    "1111100000000101",
    "1111011110110110",
    "1111011110111011",
    "1111011111111111",
    "1111100001100001",
    "1111100011001000",
    "1111100100011101",
    "1111100101001101",
    "1111100101010011",
    "1111100100101100",
    "1111100011010011",
    "1111100001001100",
    "1111011110010001",
    "1111011010100010",
    "1111010110000011",
    "1111010000111001",
    "1111001011010100",
    "1111000101100010",
    "1110111111110110",
    "1110111010100011",
    "1110110101110100",
    "1110110001110110",
    "1110101110101101",
    "1110101100010111",
    "1110101010111000",
    "1110101010000111",
    "1110101001111101",
    "1110101010001111",
    "1110101010110101",
    "1110101011101010",
    "1110101100101000",
    "1110101101110010",
    "1110101111001100",
    "1110110000111110",
    "1110110011010011",
    "1110110110001110",
    "1110111001110101",
    "1110111110000101",
    "1111000010110100",
    "1111000111111010",
    "1111001101001010",
    "1111010010010100",
    "1111010111010001",
    "1111011011111101",
    "1111100000011100",
    "1111100100110001",
    "1111101001000010",
    "1111101101010011",
    "1111110001101001",
    "1111110110000110",
    "1111111010110001",
    "1111111111110011",
    "1111111010100111",
    "1111110100011101",
    "1111101101101110",
    "1111100110101010",
    "1111011111101011",
    "1111011001001110",
    "1111010011101111",
    "1111001111011110",
    "1111001100011110",
    "1111001010100011",
    "1111001001011000",
    "1111001000101010",
    "1111001000001000",
    "1111000111100111",
    "1111000111000100",
    "1111000110100100",
    "1111000110000100",
    "1111000101100101",
    "1111000101000000",
    "1111000100001101",
    "1111000011000101",
    "1111000001011111",
    "1110111111011010",
    "1110111100111100",
    "1110111010001100",
    "1110110111011111",
    "1110110101001001",
    "1110110011100001",
    "1110110010111011",
    "1110110011100010",
    "1110110101011000",
    "1110111000011011",
    "1110111100011011",
    "1111000001001000",
    "1111000110010101",
    "1111001011110011",
    "1111010001011110",
    "1111010111010001",
    "1111011101001110",
    "1111100011010000",
    "1111101001010101",
    "1111101111010110",
    "1111110101000111",
    "1111111010011111",
    "1111111111010101",
    "1111111100011001",
    "1111111000110101",
    "1111110110000000",
    "1111110011111101",
    "1111110010101110",
    "1111110010010001",
    "1111110010100110",
    "1111110011100110",
    "1111110101001011",
    "1111110111010100",
    "1111111010000000",
    "1111111101010111",
    "1111111110011011",
    "1111111001010011",
    "1111110011000110",
    "1111101011110111",
    "1111100011101100",
    "1111011010111000",
    "1111010001110110",
    "1111001001000110",
    "1111000001001111",
    "1110111010110101",
    "1110110110010011",
    "1110110011111011",
    "1110110011100110",
    "1110110100111100",
    "1110110111100000",
    "1110111010101101",
    "1110111110000101",
    "1111000001010010",
    "1111000100001011",
    "1111000110110001",
    "1111001001000111",
    "1111001011011000",
    "1111001101100110",
    "1111001111111011",
    "1111010010010111",
    "1111010100111100",
    "1111010111101100",
    "1111011010101000",
    "1111011101101101",
    "1111100000110110",
    "1111100100000000",
    "1111100110111110",
    "1111101001101000",
    "1111101011101111",
    "1111101101000111",
    "1111101101100110",
    "1111101101000001",
    "1111101011010000",
    "1111101000001100",
    "1111100011110100",
    "1111011110000100",
    "1111010111000100",
    "1111001111000100",
    "1111000110100000",
    "1110111110000010",
    "1110110110011000",
    "1110110000010100",
    "1110101100011110",
    "1110101011010011",
    "1110101100111111",
    "1110110001011110",
    "1110111000011101",
    "1111000001011110",
    "1111001011110011",
    "1111010110101111",
    "1111100001011010",
    "1111101011000100",
    "1111110011001100",
    "1111111001100011",
    "1111111110001101",
    "1111111110100001",
    "1111111100010001",
    "1111111010101011",
    "1111111001011101",
    "1111111000100010",
    "1111110111111001",
    "1111110111101011",
    "1111110111111001",
    "1111111000100111",
    "1111111001110101",
    "1111111011100000",
    "1111111101101000",
    "1111111111110111",
    "1111111101000111",
    "1111111010001001",
    "1111110111000100",
    "1111110011111011",
    "1111110000110001",
    "1111101101100011",
    "1111101010001011",
    "1111100110100101",
    "1111100010101100",
    "1111011110011100",
    "1111011001111101",
    "1111010101010101",
    "1111010000110101",
    "1111001100101011",
    "1111001001010001",
    "1111000110110111",
    "1111000101101111",
    "1111000110000001",
    "1111000111101100",
    "1111001010100011",
    "1111001110010010",
    "1111010010100100",
    "1111010110111111",
    "1111011011001111",
    "1111011111001010",
    "1111100010100111",
    "1111100101101001",
    "1111101000010100",
    "1111101010101100",
    "1111101100110110",
    "1111101110110011",
    "1111110000100010",
    "1111110001111110",
    "1111110011000001",
    "1111110011100111",
    "1111110011101001",
    "1111110011000101",
    "1111110001111101",
    "1111110000011010",
    "1111101110100010",
    "1111101100100100",
    "1111101010101011",
    "1111101000111110",
    "1111100111100001",
    "1111100110010010",
    "1111100101001001",
    "1111100100000001",
    "1111100010110001",
    "1111100001010100",
    "1111011111110000",
    "1111011110001111",
    "1111011101000000",
    "1111011100011001",
    "1111011100101010",
    "1111011101111111",
    "1111100000011110",
    "1111100100000000",
    "1111101000010101",
    "1111101101001011",
    "1111110010001001",
    "1111110110111001",
    "1111111011000111",
    "1111111110100101",
    "1111111110110001",
    "1111111101000011",
    "1111111100000111",
    "1111111011111000",
    "1111111100001010",
    "1111111100110010",
    "1111111101101000",
    "1111111110100011",
    "1111111111011111",
    "1111111111100110",
    "1111111110110101",
    "1111111110010000",
    "1111111101111010",
    "1111111101111000",
    "1111111110001101",
    "1111111110111011",
    "1111111111110110",
    "1111111110001011",
    "1111111011111110",
    "1111111001001101",
    "1111110101110100",
    "1111110001101110",
    "1111101100110111",
    "1111100111001101",
    "1111100000101011",
    "1111011001010101",
    "1111010001001111",
    "1111001000100011",
    "1110111111100001",
    "1110110110010110",
    "1110101101010110",
    "1110100100110011",
    "1110011100111000",
    "1110010101110100",
    "1110001111101001",
    "1110001010011101",
    "1110000110001110",
    "1110000011000001",
    "1110000000110101",
    "1101111111101000",
    "1101111111010100",
    "1101111111110001",
    "1110000000110011",
    "1110000010000101",
    "1110000011011100",
    "1110000100101100",
    "1110000101101111",
    "1110000110101000",
    "1110000111100010",
    "1110001000101000",
    "1110001010000100",
    "1110001100000100",
    "1110001110110000",
    "1110010010001101",
    "1110010110100000",
    "1110011011110000",
    "1110100010000010",
    "1110101001010110",
    "1110110001101100",
    "1110111010110010",
    "1111000100010011",
    "1111001101101101",
    "1111010110100000",
    "1111011110001010",
    "1111100100010011",
    "1111101000110001",
    "1111101011100101",
    "1111101100111111",
    "1111101101011010",
    "1111101101001110",
    "1111101100110101",
    "1111101100100000",
    "1111101100011011",
    "1111101100101001",
    "1111101101001101",
    "1111101110000110",
    "1111101111010110",
    "1111110000111010",
    "1111110010110011",
    "1111110100111001",
    "1111110111000100",
    "1111111001001001",
    "1111111010111101",
    "1111111100010111",
    "1111111101011001",
    "1111111110000110",
    "1111111110101101",
    "1111111111100000",
    "1111111111001111",
    "1111111101011010",
    "1111111010111110",
    "1111111000000100",
    "1111110100111111",
    "1111110010001010",
    "1111101111111010",
    "1111101110100001",
    "1111101110000110",
    "1111101110100111",
    "1111101111111001",
    "1111110001110010",
    "1111110100000111",
    "1111110110110011",
    "1111111001110010",
    "1111111101000100",
    "1111111111011000",
    "1111111011101100",
    "1111110111111110",
    "1111110100011010",
    "1111110001001110",
    "1111101110101000",
    "1111101100101111",
    "1111101011101010",
    "1111101011011100",
    "1111101100000011",
    "1111101101011100",
    "1111101111011110",
    "1111110001111100",
    "1111110100100110",
    "1111110111001000",
    "1111111001010101",
    "1111111011000001",
    "1111111100001000",
    "1111111100101110",
    "1111111101000011",
    "1111111101010110",
    "1111111101111000",
    "1111111110110110",
    "1111111111101000",
    "1111111101110001",
    "1111111011110000",
    "1111111001111001",
    "1111111000100101",
    "1111111000001000",
    "1111111000110011",
    "1111111010110011",
    "1111111110001110",
    "1111111100110001",
    "1111110110001110",
    "1111101110001111",
    "1111100101000101",
    "1111011011001100",
    "1111010001001100",
    "1111000111101100",
    "1110111111001010",
    "1110110111111010",
    "1110110001111011",
    "1110101101000000",
    "1110101000111100",
    "1110100101011111",
    "1110100010100111",
    "1110100000011010",
    "1110011111000010",
    "1110011110101000",
    "1110011111001100",
    "1110100000101110",
    "1110100011000101",
    "1110100110000011",
    "1110101001100000",
    "1110101101011001",
    "1110110001100110",
    "1110110110000110",
    "1110111010110010",
    "1110111111100001",
    "1111000100001000",
    "1111001000011110",
    "1111001100011011",
    "1111001111110101",
    "1111010010101110",
    "1111010101000101",
    "1111010110111111",
    "1111011000100111",
    "1111011001111111",
    "1111011011010100",
    "1111011100101010",
    "1111011110000010",
    "1111011111100001",
    "1111100001000101",
    "1111100010110100",
    "1111100100110100",
    "1111100111001000",
    "1111101001111101",
    "1111101101011001",
    "1111110001011011",
    "1111110101111110",
    "1111111010110100",
    "1111111111101000",
    "1111111011111001",
    "1111111000001001",
    "1111110101010011",
    "1111110011011010",
    "1111110010010100",
    "1111110001110010",
    "1111110001011101",
    "1111110000111111",
    "1111110000000100",
    "1111101110011111",
    "1111101100001010",
    "1111101001000010",
    "1111100101010000",
    "1111100000111101",
    "1111011100010100",
    "1111010111100000",
    "1111010010101110",
    "1111001101111101",
    "1111001001010011",
    "1111000100100111",
    "1110111111110101",
    "1110111010110101",
    "1110110101101010",
    "1110110000100001",
    "1110101011110010",
    "1110100111111111",
    "1110100101101010",
    "1110100101010011",
    "1110100111001110",
    "1110101011011001",
    "1110110001100100",
    "1110111001001001",
    "1111000001011100",
    "1111001001100111",
    "1111010000111000",
    "1111010110100111",
    "1111011010011110",
    "1111011100011011",
    "1111011100101000",
    "1111011011100011",
    "1111011001100101",
    "1111010111001001",
    "1111010100100100",
    "1111010001111101",
    "1111001111010100",
    "1111001100100110",
    "1111001001110010",
    "1111000110110010",
    "1111000011100100",
    "1111000000001010",
    "1110111100100110",
    "1110111000111111",
    "1110110101011011",
    "1110110010000011",
    "1110101111000010",
    "1110101100100110",
    "1110101010111100",
    "1110101010001001",
    "1110101010001111",
    "1110101011001110",
    "1110101100111000",
    "1110101111001000",
    "1110110001111000",
    "1110110101000001",
    "1110111000100010",
    "1110111100011100",
    "1111000000110000",
    "1111000101010011",
    "1111001001111101",
    "1111001110011110",
    "1111010010100001",
    "1111010101110111",
    "1111011000010011",
    "1111011001101101",
    "1111011010000111",
    "1111011001101011",
    "1111011000100101",
    "1111010110111111",
    "1111010101000101",
    "1111010010111101",
    "1111010000101110",
    "1111001110011111",
    "1111001100010011",
    "1111001010001100",
    "1111001000010001",
    "1111000110100000",
    "1111000100110100",
    "1111000011000101",
    "1111000001001101",
    "1110111111001000",
    "1110111100110101",
    "1110111010011101",
    "1110111000010000",
    "1110110110100000",
    "1110110101100000",
    "1110110101011101",
    "1110110110011111",
    "1110111000011110",
    "1110111011010100",
    "1110111110101011",
    "1111000010010100",
    "1111000101111100",
    "1111001001011110",
    "1111001100110111",
    "1111010000010001",
    "1111010011111000",
    "1111010111111100",
    "1111011100101000",
    "1111100001111110",
    "1111100111111001",
    "1111101110001011",
    "1111110100100000",
    "1111111010100111",
    "1111111111110000",
    "1111111010110101",
    "1111110110101110",
    "1111110011011011",
    "1111110000111011",
    "1111101111001100",
    "1111101110000111",
    "1111101101101010",
    "1111101101110001",
    "1111101110011101",
    "1111101111110000",
    "1111110001110101",
    "1111110100111100",
    "1111111001010101",
    "1111111111010101",
    "1111111000111010",
    "1111101111101010",
    "1111100101011101",
    "1111011011010100",
    "1111010010010010",
    "1111001011011000",
    "1111000111001000",
    "1111000101100000",
    "1111000110000001",
    "1111000111110010",
    "1111001001111101",
    "1111001011111100",
    "1111001101011011",
    "1111001110011111",
    "1111001111011001",
    "1111010000011010",
    "1111010001110001",
    "1111010011011101",
    "1111010101011010",
    "1111010111011010",
    "1111011001010000",
    "1111011010101111",
    "1111011011110010",
    "1111011100011001",
    "1111011100101010",
    "1111011100110000",
    "1111011100111101",
    "1111011101100110",
    "1111011111000000",
    "1111100001011110",
    "1111100101001011",
    "1111101010001110",
    "1111110000100000",
    "1111110111110011",
    "1111111111101110",
    "1111111000000111",
    "1111110000010010",
    "1111101001001101",
    "1111100011001011",
    "1111011110010010",
    "1111011010100000",
    "1111010111100000",
    "1111010101000000",
    "1111010010100111",
    "1111010000001010",
    "1111001101100011",
    "1111001010111000",
    "1111001000011101",
    "1111000110100000",
    "1111000101010101",
    "1111000101001000",
    "1111000110000001",
    "1111000111111100",
    "1111001010110100",
    "1111001110100001",
    "1111010010111001",
    "1111010111110010",
    "1111011101000100",
    "1111100010100111",
    "1111101000010000",
    "1111101101110100",
    "1111110011000110",
    "1111110111111010",
    "1111111100001101",
    "1111111111111011",
    "1111111100110101",
    "1111111010000111",
    "1111110111110111",
    "1111110110000100",
    "1111110100110101",
    "1111110100001101",
    "1111110100010000",
    "1111110100111011",
    "1111110110001010",
    "1111110111110101",
    "1111111001111010",
    "1111111100010100",
    "1111111111000110",
    "1111111101100111",
    "1111111001101100",
    "1111110100111100",
    "1111101111001101",
    "1111101000010101",
    "1111100000010101",
    "1111010111010101",
    "1111001101100100",
    "1111000011100010",
    "1110111001110111",
    "1110110001001100",
    "1110101010000111",
    "1110100101000110",
    "1110100010010010",
    "1110100001100111",
    "1110100010110110",
    "1110100101100010",
    "1110101001010000",
    "1110101101100011",
    "1110110010000000",
    "1110110110010000",
    "1110111010000010",
    "1110111101001001",
    "1110111111011010",
    "1111000000101110",
    "1111000001000101",
    "1111000000011001",
    "1110111110101000",
    "1110111011110010",
    "1110110111111010",
    "1110110011001101",
    "1110101101111011",
    "1110101000100011",
    "1110100011100100",
    "1110011111011100",
    "1110011100100001",
    "1110011011000100",
    "1110011011000110",
    "1110011100100001",
    "1110011111001000",
    "1110100010101111",
    "1110100111001000",
    "1110101100000100",
    "1110110001010100",
    "1110110110101010",
    "1110111011110010",
    "1111000000010101",
    "1111000100000011",
    "1111000110101101",
    "1111001000010000",
    "1111001000110100",
    "1111001000101100",
    "1111001000010001",
    "1111001000000110",
    "1111001000100010",
    "1111001001111010",
    "1111001100010100",
    "1111001111110001",
    "1111010100000101",
    "1111011001000001",
    "1111011110010111",
    "1111100100000000",
    "1111101001110000",
    "1111101111100111",
    "1111110101100011",
    "1111111011011100",
    "1111111110110110",
    "1111111001101011",
    "1111110101010001",
    "1111110001110100",
    "1111101111011000",
    "1111101101110111",
    "1111101100111101",
    "1111101100011001",
    "1111101011110111",
    "1111101011001010",
    "1111101010001101",
    "1111101000111110",
    "1111100111100000",
    "1111100101110100",
    "1111100011111001",
    "1111100001110001",
    "1111011111011010",
    "1111011100110101",
    "1111011010000111",
    "1111010111011000",
    "1111010100101110",
    "1111010010010000",
    "1111010000000101",
    "1111001110001111",
    "1111001100110011",
    "1111001011110010",
    "1111001011001010",
    "1111001010111101",
    "1111001011001010",
    "1111001011110010",
    "1111001100111000",
    "1111001110011100",
    "1111010000100001",
    "1111010011000101",
    "1111010110000100",
    "1111011001011110",
    "1111011101001010",
    "1111100000111110",
    "1111100100110001",
    "1111101000011001",
    "1111101011101101",
    "1111101110101001",
    "1111110001001101",
    "1111110011011110",
    "1111110101100101",
    "1111110111101011",
    "1111111001111001",
    "1111111100010001",
    "1111111110110110",
    "1111111110011011",
    "1111111011101110",
    "1111111001001010",
    "1111110110110100",
    "1111110100110110",
    "1111110011010001",
    "1111110010000110",
    "1111110001001110",
    "1111110000100010",
    "1111101111110101",
    "1111101110111010",
    "1111101101100100",
    "1111101011101001",
    "1111101001000011",
    "1111100101110010",
    "1111100001111011",
    "1111011101100001",
    "1111011000110100",
    "1111010011111000",
    "1111001110110101",
    "1111001001101111",
    "1111000100100111",
    "1110111111011110",
    "1110111010010100",
    "1110110101010000",
    "1110110000010100",
    "1110101011110000",
    "1110100111101100",
    "1110100100010101",
    "1110100001110001",
    "1110100000000010",
    "1110011111000111",
    "1110011110111000",
    "1110011111010001",
    "1110100000001010",
    "1110100001100110",
    "1110100011100111",
    "1110100110001011",
    "1110101001011000",
    "1110101101000111",
    "1110110001010100",
    "1110110101110110",
    "1110111010100000",
    "1110111111000111",
    "1111000011100110",
    "1111000111110111",
    "1111001011111111",
    "1111010000000111",
    "1111010100011010",
    "1111011001000110",
    "1111011110011011",
    "1111100100011111",
    "1111101011011100",
    "1111110011001110",
    "1111111011101010",
    "1111111011100011",
    "1111110011000000",
    "1111101011001111",
    "1111100100101111",
    "1111011111110110",
    "1111011100101011",
    "1111011011000010",
    "1111011010101000",
    "1111011010111101",
    "1111011011101010",
    "1111011100010110",
    "1111011100110000",
    "1111011100101101",
    "1111011100000010",
    "1111011010101101",
    "1111011000101111",
    "1111010110001000",
    "1111010011000000",
    "1111001111100011",
    "1111001011111010",
    "1111001000010000",
    "1111000100100100",
    "1111000000101110",
    "1110111100100001",
    "1110110111110010",
    "1110110010100001",
    "1110101100111111",
    "1110100111110101",
    "1110100011111100",
    "1110100010010000",
    "1110100011100111",
    "1110101000100111",
    "1110110001011001",
    "1110111101100001",
    "1111001011111010",
    "1111011011000010",
    "1111101001001011",
    "1111110100110110",
    "1111111101010001",
    "1111111101100110",
    "1111111011000111",
    "1111111010000110",
    "1111111001011011",
    "1111111000010100",
    "1111110110100001",
    "1111110100010011",
    "1111110010001000",
    "1111110000100011",
    "1111101111111001",
    "1111110000001111",
    "1111110001011000",
    "1111110011000110",
    "1111110101000110",
    "1111110111010001",
    "1111111001101000",
    "1111111100010111",
    "1111111111101011",
    "1111111100000111",
    "1111110110110111",
    "1111110000011001",
    "1111101000110001",
    "1111100000010010",
    "1111010111100000",
    "1111001111001111",
    "1111001000011011",
    "1111000100000000",
    "1111000010100001",
    "1111000100001000",
    "1111001000010110",
    "1111001110010110",
    "1111010101000001",
    "1111011011011110",
    "1111100001000111",
    "1111100101101010",
    "1111101001001110",
    "1111101011111000",
    "1111101101101101",
    "1111101110100111",
    "1111101110011101",
    "1111101101000111",
    "1111101010100101",
    "1111100110111110",
    "1111100010100110",
    "1111011101110010",
    "1111011000111111",
    "1111010100101100",
    "1111010001001100",
    "1111001110100100",
    "1111001100110011",
    "1111001011100011",
    "1111001010011000",
    "1111001000110101",
    "1111000110101111",
    "1111000100000101",
    "1111000001000011",
    "1110111110001001",
    "1110111011101000",
    "1110111001110010",
    "1110111000101000",
    "1110111000000011",
    "1110110111111001",
    "1110111000001000",
    "1110111001000010",
    "1110111011011000",
    "1111000000000011",
    "1111000111111001",
    "1111010011000001",
    "1111100000101100",
    "1111101111010101",
    "1111111101000000",
    "1111110111111001",
    "1111110000011010",
    "1111101100100011",
    "1111101100000101",
    "1111101111001110",
    "1111110111000100",
    "1111111011000110",
    "1111100111000100",
    "1111001110100011",
    "1110110101011000",
    "1110100000011111",
    "1110010100011010",
    "1110010011101100",
    "1110011110001001",
    "1110110001000101",
    "1111001000100101",
    "1111100000101011",
    "1111110110001101",
    "1111111000100111",
    "1111101100101110",
    "1111100110001101",
    "1111100100101111",
    "1111100111110011",
    "1111101110011101",
    "1111110111100001",
    "1111111110011010",
    "1111110101000100",
    "1111101101110101",
    "1111101001101000",
    "1111101000100010",
    "1111101001111001",
    "1111101100100100",
    "1111101111010000",
    "1111110000100110",
    "1111101111010111",
    "1111101010110010",
    "1111100011000000",
    "1111011001001110",
    "1111001111010111",
    "1111000111100010",
    "1111000011010111",
    "1111000011010000",
    "1111000110100000",
    "1111001011011011",
    "1111010000001010",
    "1111010011011100",
    "1111010101000000",
    "1111010101100100",
    "1111010110010110",
    "1111011000101101",
    "1111011101010110",
    "1111100100000011",
    "1111101011110110",
    "1111110011010010",
    "1111111001000100",
    "1111111100100010",
    "1111111101101011",
    "1111111100111110",
    "1111111011000110",
    "1111111000101011",
    "1111110110001000",
    "1111110011101010",
    "1111110001001100",
    "1111101110011010",
    "1111101010111101",
    "1111100110100111",
    "1111100001011111",
    "1111011011111111",
    "1111010110110010",
    "1111010010100100",
    "1111001111101110",
    "1111001110011100",
    "1111001110011111",
    "1111001111101000",
    "1111010001100010",
    "1111010100001110",
    "1111010111111010",
    "1111011100110011",
    "1111100010111110",
    "1111101010001101",
    "1111110001111100",
    "1111111001010101",
    "1111111111010110",
    "1111111101000010",
    "1111111100101010",
    "1111111111110111",
    "1111111001100100",
    "1111110000100101",
    "1111100110101001",
    "1111011101100011",
    "1111010111000011",
    "1111010100010000",
    "1111010101011111",
    "1111011010000111",
    "1111100000110110",
    "1111101000000010",
    "1111101110000111",
    "1111110010000001",
    "1111110011011111",
    "1111110010111001",
    "1111110001000101",
    "1111101110111111",
    "1111101101011011",
    "1111101100110111",
    "1111101101111010",
    "1111110010000110",
    "1111111100000101",
    "1111110001101011",
    "1111010110101100",
    "1110110101010101",
    "1110010010100111",
    "1101110100011111",
    "1101100000000010",
    "1101010111101100",
    "1101011010100011",
    "1101100101110001",
    "1101110110100010",
    "1110001011001001",
    "1110100010110001",
    "1110111100010111",
    "1111010101110001",
    "1111101011101011",
    "1111111010100010",
    "1111111111110000",
    "1111111011001001",
    "1111101111010010",
    "1111100000010010",
    "1111010010011100",
    "1111001000100000",
    "1111000010110011",
    "1110111111011010",
    "1110111011010001",
    "1110110011101001",
    "1110100111110111",
    "1110011001101000",
    "1110001100010001",
    "1110000011100110",
    "1110000010100010",
    "1110001010010001",
    "1110011001111010",
    "1110101110110101",
    "1111000101011011",
    "1111011010000001",
    "1111101001010111",
    "1111110001010010",
    "1111110000110000",
    "1111100111111101",
    "1111011000001001",
    "1111000011100001",
    "1110101100111100",
    "1110010111101000",
    "1110000110100111",
    "1101111011111101",
    "1101111000100010",
    "1101111011111101",
    "1110000100110100",
    "1110010001001111",
    "1110011111011100",
    "1110101101111010",
    "1110111011100000",
    "1111000111011111",
    "1111010001010111",
    "1111011001000110",
    "1111011110111011",
    "1111100011011101",
    "1111100111010010",
    "1111101010110101",
    "1111101110001101",
    "1111110001001101",
    "1111110011011110",
    "1111110100101110",
    "1111110100110101",
    "1111110011110001",
    "1111110001101001",
    "1111101110100000",
    "1111101010011111",
    "1111100101101001",
    "1111100000010100",
    "1111011011010001",
    "1111010111001001",
    "1111010100001101",
    "1111010001111011",
    "1111001111010010",
    "1111001011001001",
    "1111000100100100",
    "1110111011010011",
    "1110101111110000",
    "1110100010111110",
    "1110010110001000",
    "1110001010100010",
    "1110000001100010",
    "1101111100110010",
    "1101111110000100",
    "1110000110110110",
    "1110011000000001",
    "1110110001011010",
    "1111010001010111",
    "1111110100011001",
    "1111101010000010",
    "1111001110100110",
    "1110111100100000",
    "1110110100101100",
    "1110110101110100",
    "1110111100110101",
    "1111000110000000",
    "1111001110001111",
    "1111010011110001",
    "1111010110010110",
    "1111010110101000",
    "1111010110110001",
    "1111011010110111",
    "1111100111010011",
    "1111111101111011",
    "1111100011000110",
    "1111000001011111",
    "1110100100011010",
    "1110010010010100",
    "1110001110111000",
    "1110011001000110",
    "1110101011110010",
    "1111000000001010",
    "1111010000010111",
    "1111011001000111",
    "1111011010010110",
    "1111010110000000",
    "1111001110111010",
    "1111000111101010",
    "1111000001010111",
    "1110111011111101",
    "1110110111000110",
    "1110110010011010",
    "1110101110011100",
    "1110101100010011",
    "1110101100111010",
    "1110110010001111",
    "1111000000000111",
    "1111011001010001",
    "1111111101100000",
    "1111010111100101",
    "1110101110010110",
    "1110001111100001",
    "1110000010010101",
    "1110001010111010",
    "1110100111010011",
    "1111010000001000",
    "1111111011100101",
    "1111100000000101",
    "1111001001001011",
    "1111000001010100",
    "1111000110100000",
    "1111010011010111",
    "1111100001010100",
    "1111101011101111",
    "1111110010010011",
    "1111111001111100",
    "1111110111001000",
    "1111011110010001",
    "1110111101101000",
    "1110011011101101",
    "1110000000000111",
    "1101110000111011",
    "1101110000100100",
    "1101111100101000",
    "1110001111011111",
    "1110100011010111",
    "1110110011111011",
    "1110111111010100",
    "1111000100101111",
    "1111000011101100",
    "1110111100001001",
    "1110101110110110",
    "1110011101101001",
    "1110001011100011",
    "1101111011110000",
    "1101110000100110",
    "1101101010110100",
    "1101101001011000",
    "1101101010010011",
    "1101101011100001",
    "1101101100001100",
    "1101101101001001",
    "1101110000001000",
    "1101110110010110",
    "1110000000101100",
    "1110010001111110",
    "1110101100111010",
    "1111010001101001",
    "1111111101001110",
    "1111010110110001",
    "1110110001110100",
    "1110011001110010",
    "1110010010001011",
    "1110011001111100",
    "1110101011100001",
    "1111000000000101",
    "1111010001101100",
    "1111011101010111",
    "1111100100011100",
    "1111101100000100",
    "1111111011000111",
    "1111101010010000",
    "1111000101010010",
    "1110011100000001",
    "1101110111001110",
    "1101011111000100",
    "1101011000010011",
    "1101100001110001",
    "1101110101000001",
    "1110001010011011",
    "1110011100010100",
    "1110101000101100",
    "1110110000101001",
    "1110110101110001",
    "1110111001001011",
    "1110111010110111",
    "1110111001001110",
    "1110110010110110",
    "1110100111111110",
    "1110011010111100",
    "1110001111101100",
    "1110001001111101",
    "1110001011011011",
    "1110010011010111",
    "1110011111011001",
    "1110101101000111",
    "1110111010111000",
    "1111000111101101",
    "1111010010101110",
    "1111011011000010",
    "1111011111111011",
    "1111100001001101",
    "1111011111101000",
    "1111011100100000",
    "1111011001001001",
    "1111010110010110",
    "1111010100011100",
    "1111010011000000",
    "1111010001101100",
    "1111010000011010",
    "1111001111101001",
    "1111001111111111",
    "1111010010101111",
    "1111011010111100",
    "1111101011100110",
    "1111111010101111",
    "1111011010110101",
    "1110111010000001",
    "1110011110001111",
    "1110001011111000",
    "1110000100101010",
    "1110000110101010",
    "1110001100111100",
    "1110010010100010",
    "1110010100010010",
    "1110010010001101",
    "1110010000111110",
    "1110010111000011",
    "1110101000011010",
    "1111000100011100",
    "1111100101011111",
    "1111111100100010",
    "1111101000101101",
    "1111100011000101",
    "1111101010101111",
    "1111111010011001",
    "1111110011011000",
    "1111100001000011",
    "1111001101111010",
    "1110111000001011",
    "1110100000001000",
    "1110001000100101",
    "1101110101100100",
    "1101101011100101",
    "1101101101011110",
    "1101111010011011",
    "1110001110110011",
    "1110100101011000",
    "1110111001001011",
    "1111000111110101",
    "1111010001110100",
    "1111011001011011",
    "1111100001111011",
    "1111101110010010",
    "1111111111101010",
    "1111101010111000",
    "1111010100101111",
    "1111000010001010",
    "1110110110101101",
    "1110110100101010",
    "1110111100001010",
    "1111001011001110",
    "1111011110010010",
    "1111110001011110",
    "1111111110110001",
    "1111110100011110",
    "1111110000000001",
    "1111110000100111",
    "1111110100110001",
    "1111111010111000",
    "1111111111111110",
    "1111111111101100",
    "1111110110110000",
    "1111100100100100",
    "1111001011110000",
    "1110110001001010",
    "1110011010000111",
    "1110001011001100",
    "1110000110100101",
    "1110001010101101",
    "1110010011101001",
    "1110011101001111",
    "1110100100100100",
    "1110101000101101",
    "1110101010001011",
    "1110101001101000",
    "1110100111111110",
    "1110100101011111",
    "1110100010001101",
    "1110011110010001",
    "1110011010001001",
    "1110010110111110",
    "1110010111100101",
    "1110011111111010",
    "1110110010011001",
    "1111001110001001",
    "1111101110110011",
    "1111110010001001",
    "1111011011101011",
    "1111010011010010",
    "1111011010110010",
    "1111101110101100",
    "1111111000110011",
    "1111100101010000",
    "1111011110011110",
    "1111101000000100",
    "1111111110111111",
    "1111011011110111",
    "1110110110010101",
    "1110010110001000",
    "1110000000011111",
    "1101110111001110",
    "1101111000111010",
    "1110000010010101",
    "1110001111011111",
    "1110011100110010",
    "1110100111010011",
    "1110101111000010",
    "1110110111101010",
    "1111000101001011",
    "1111011001010101",
    "1111110010011001",
    "1111110101000000",
    "1111100100101110",
    "1111100100101110",
    "1111111001001111",
    "1111100000100110",
    "1110110001111101",
    "1110000110010011",
    "1101100111101101",
    "1101011011000111",
    "1101011111011111",
    "1101110000011111",
    "1110001001110111",
    "1110101000010110",
    "1111001001111101",
    "1111101101001001",
    "1111110000010000",
    "1111010001000011",
    "1110111000100000",
    "1110101001011101",
    "1110100011110011",
    "1110100100100111",
    "1110101000001000",
    "1110101011010011",
    "1110101100111100",
    "1110101101011100",
    "1110101110111011",
    "1110110101100100",
    "1111000100101100",
    "1111011100010011",
    "1111111000100010",
    "1111101101110001",
    "1111011110101110",
    "1111011111101100",
    "1111110001010010",
    "1111110001001101",
    "1111010000000010",
    "1110110011100110",
    "1110100010010100",
    "1110011110000111",
    "1110100100000001",
    "1110101110011111",
    "1110111000001011",
    "1110111110000010",
    "1111000000010101",
    "1111000001011111",
    "1111000100011010",
    "1111001011001110",
    "1111010101110110",
    "1111100010000011",
    "1111101100111101",
    "1111110100001011",
    "1111110110110100",
    "1111110101011000",
    "1111110001000010",
    "1111101011100000",
    "1111100110101111",
    "1111100011111000",
    "1111100011000000",
    "1111100011010000",
    "1111100011011101",
    "1111100101001001",
    "1111101100101100",
    "1111111101110111",
    "1111100110001000",
    "1111000010000101",
    "1110011011111101",
    "1101111010101011",
    "1101100100001010",
    "1101011011001010",
    "1101011101110011",
    "1101100111011101",
    "1101110011001010",
    "1101111101010110",
    "1110000101010101",
    "1110001011101101",
    "1110010001011100",
    "1110010111100011",
    "1110011110000101",
    "1110100100000000",
    "1110100111011101",
    "1110100111111111",
    "1110101001010001",
    "1110110000010010",
    "1110111111111000",
    "1111010111010101",
    "1111110001110011",
    "1111110110101001",
    "1111100110101011",
    "1111100000100100",
    "1111100010001111",
    "1111100110101000",
    "1111101000111101",
    "1111100110000000",
    "1111011101101001",
    "1111010010000101",
    "1111000110010000",
    "1111000000001111",
    "1111000101111001",
    "1111011000110101",
    "1111110110110110",
    "1111100110000011",
    "1111000101100101",
    "1110101101100110",
    "1110100001100110",
    "1110100001000011",
    "1110101000000001",
    "1110110001111001",
    "1110111010011000",
    "1110111110011110",
    "1110111110001010",
    "1110111010100110",
    "1110110101110001",
    "1110110001100010",
    "1110101110000100",
    "1110101010010001",
    "1110100101000011",
    "1110011101101011",
    "1110010100011101",
    "1110001011000100",
    "1110000011101100",
    "1110000000000010",
    "1110000000110001",
    "1110000101100101",
    "1110001101010010",
    "1110011000010001",
    "1110101000111010",
    "1111000000111000",
    "1111011111111010",
    "1111111100111001",
    "1111011010101010",
    "1110111110011100",
    "1110101100100001",
    "1110100110101010",
    "1110101010000110",
    "1110110001111101",
    "1110111001110100",
    "1110111110101001",
    "1111000000011110",
    "1111000000011110",
    "1111000000001111",
    "1111000100101110",
    "1111010010010101",
    "1111101001110011",
    "1111110111100101",
    "1111011000100010",
    "1111000000110001",
    "1110110101110010",
    "1110111100001111",
    "1111010110011010",
    "1111111110100000",
    "1111001001100101",
    "1110010100110011",
    "1101101011111100",
    "1101011001100101",
    "1101100100010011",
    "1110001010110111",
    "1111000010101110",
    "1111111101000101",
    "1111010011100010",
    "1110111000001011",
    "1110110010010101",
    "1110111100101010",
    "1111001110110011",
    "1111100000100011",
    "1111101100010111",
    "1111110001100010",
    "1111110010100001",
    "1111110010100111",
    "1111110111001000",
    "1111111011000101",
    "1111100011000011",
    "1111000010101011",
    "1110011110101101",
    "1101111101101000",
    "1101100101010010",
    "1101011010001011",
    "1101011101010110",
    "1101101011001100",
    "1101111110010001",
    "1110010000110101",
    "1110011110101000",
    "1110100110110001",
    "1110101010010001",
    "1110101010110010",
    "1110101010100101",
    "1110101010100010",
    "1110101010110000",
    "1110101101000101",
    "1110110011111011",
    "1111000000010111",
    "1111010001100100",
    "1111100100011101",
    "1111110101000011",
    "1111111111100011",
    "1111111010010011",
    "1111111000101111",
    "1111110110000101",
    "1111101110110011",
    "1111100001110100",
    "1111010001010100",
    "1111000001101110",
    "1110110111000011",
    "1110110011011111",
    "1110110110101101",
    "1110111101101001",
    "1111000100100010",
    "1111001000101000",
    "1111001000101010",
    "1111000101101100",
    "1111000010000010",
    "1111000001010010",
    "1111001001000100",
    "1111011101010110",
    "1111111110000100",
    "1111011000011000",
    "1110101101100001",
    "1110001001100011",
    "1101110011001010",
    "1101101101111000",
    "1101110111101000",
    "1110001001110101",
    "1110011101000000",
    "1110101010011110",
    "1110101110100110",
    "1110101001111010",
    "1110011110101101",
    "1110010001000011",
    "1110000111110101",
    "1110001001111100",
    "1110011010111000",
    "1110111001101000",
    "1111011111111000",
    "1111111010111101",
    "1111011110010010",
    "1111001111001000",
    "1111001110001111",
    "1111010111001101",
    "1111100011100001",
    "1111101100110111",
    "1111101111101111",
    "1111101100011000",
    "1111100100100101",
    "1111011010101011",
    "1111010001000101",
    "1111001000011101",
    "1111000000100001",
    "1110111001001011",
    "1110110010010010",
    "1110101100100001",
    "1110101001001011",
    "1110101001000111",
    "1110101100010111",
    "1110110001011010",
    "1110110111001101",
    "1111000000001101",
    "1111010000011001",
    "1111101001101111",
    "1111110100011010",
    "1111001110011100",
    "1110101010101101",
    "1110001111011010",
    "1110000001100001",
    "1110000001100010",
    "1110001011001110",
    "1110011000101111",
    "1110100100101111",
    "1110101100100011",
    "1110110000111110",
    "1110110011110110",
    "1110110111011010",
    "1110111101011011",
    "1111000101100101",
    "1111001110000000",
    "1111010100011111",
    "1111010111001110",
    "1111010110000011",
    "1111010010000110",
    "1111001100101101",
    "1111000110101100",
    "1111000000100011",
    "1110111011000001",
    "1110110111001110",
    "1110110110000001",
    "1110110111101111",
    "1110111011110111",
    "1111000010111011",
    "1111010000000111",
    "1111100110001101",
    "1111111011000000",
    "1111010110111001",
    "1110110011101111",
    "1110011000100000",
    "1110001010110000",
    "1110001101001010",
    "1110011100100000",
    "1110110001101100",
    "1111000101111001",
    "1111010011111011",
    "1111011010001110",
    "1111011010010011",
    "1111010110111011",
    "1111010011010111",
    "1111010001111011",
    "1111010010010101",
    "1111010011000110",
    "1111010010010111",
    "1111001110110001",
    "1111001000011101",
    "1111000000101011",
    "1110111000110101",
    "1110110001101001",
    "1110101100111010",
    "1110101111000101",
    "1110111100001001",
    "1111010100100111",
    "1111110100111111",
    "1111101001010101",
    "1111001101100100",
    "1110111101000111",
    "1110111010110000",
    "1111000101100000",
    "1111011000001100",
    "1111101011010011",
    "1111110111101001",
    "1111111001011100",
    "1111110001000110",
    "1111100010001101",
    "1111010010001101",
    "1111000110101111",
    "1111000010111011",
    "1111000101111100",
    "1111001100000010",
    "1111010000101001",
    "1111010000111101",
    "1111001111001111",
    "1111010001011110",
    "1111011100010011",
    "1111110001101111",
    "1111110000010010",
    "1111001111101001",
    "1110110010111000",
    "1110011111111000",
    "1110011001010011",
    "1110011100001111",
    "1110100011000101",
    "1110101000101111",
    "1110101010011011",
    "1110101010001100",
    "1110101101111011",
    "1110111010111100",
    "1111010011101010",
    "1111110101100101",
    "1111100110101000",
    "1111001000110101",
    "1110110111010110",
    "1110110100111011",
    "1110111110100110",
    "1111010000101011",
    "1111101001111101",
    "1111110110001101",
    "1111010000110110",
    "1110101000111100",
    "1110000100101100",
    "1101101001111001",
    "1101011101100011",
    "1101100001111101",
    "1101110011011100",
    "1110001011001110",
    "1110100010001011",
    "1110110010110100",
    "1110111011101111",
    "1110111110010010",
    "1110111101010110",
    "1110111100011001",
    "1110111101010100",
    "1110111111110110",
    "1111000011000000",
    "1111000101011011",
    "1111000110100101",
    "1111000111011000",
    "1111001001110101",
    "1111010001001100",
    "1111100000000011",
    "1111110110101000",
    "1111101101000100",
    "1111001111000111",
    "1110110100010000",
    "1110100000010010",
    "1110010101000011",
    "1110010000111011",
    "1110010000110101",
    "1110010100000110",
    "1110011100001110",
    "1110101010100110",
    "1110111110101110",
    "1111010100001011",
    "1111100101010010",
    "1111101110110010",
    "1111110000110001",
    "1111110000000001",
    "1111110100001110",
    "1111111101001000",
    "1111100011011100",
    "1111000011011000",
    "1110100101101111",
    "1110010010010010",
    "1110001101000100",
    "1110010100111011",
    "1110100011100001",
    "1110110001001010",
    "1110111000011010",
    "1110110111000011",
    "1110101110110001",
    "1110100100000001",
    "1110011010110000",
    "1110010101001110",
    "1110010110001101",
    "1110100000101011",
    "1110110110001000",
    "1111010101101010",
    "1111111011001010",
    "1111011111011110",
    "1111000000001010",
    "1110101011100101",
    "1110100010101110",
    "1110100010010101",
    "1110100101011000",
    "1110100111000011",
    "1110100100011101",
    "1110011101110000",
    "1110010100101010",
    "1110001011110101",
    "1110000110001101",
    "1110000100101110",
    "1110000110110111",
    "1110001101110111",
    "1110011100011011",
    "1110110100100010",
    "1111010110001000",
    "1111111101011111",
    "1111011100010111",
    "1110111111000111",
    "1110110000110001",
    "1110110010110110",
    "1111000000101110",
    "1111010011001101",
    "1111100011010111",
    "1111101100100111",
    "1111101110110011",
    "1111101011101001",
    "1111100110111100",
    "1111100111110110",
    "1111110011100011",
    "1111110101001110",
    "1111010101100101",
    "1110110100010010",
    "1110010111110111",
    "1110000100111011",
    "1101111101010100",
    "1110000000000011",
    "1110001100110010",
    "1110100011100001",
    "1111000001110100",
    "1111100011111001",
    "1111111011011101",
    "1111100001110110",
    "1111010010011111",
    "1111001110001111",
    "1111010010111001",
    "1111011011100000",
    "1111100011110001",
    "1111101000111111",
    "1111101010100101",
    "1111101100010100",
    "1111110100000001",
    "1111111010001000",
    "1111011101111111",
    "1110111101000100",
    "1110011111110110",
    "1110001101010001",
    "1110001001011000",
    "1110010011010010",
    "1110100100111011",
    "1110110111100111",
    "1111000110110010",
    "1111010000111011",
    "1111010111000100",
    "1111011011110111",
    "1111100100101010",
    "1111110111001010",
    "1111101011101010",
    "1111000111101010",
    "1110100100100010",
    "1110001011000001",
    "1110000001000010",
    "1110001000010110",
    "1110011101000010",
    "1110110111000110",
    "1111001110111000",
    "1111011110010110",
    "1111100010101110",
    "1111011100111000",
    "1111001111100011",
    "1110111110111010",
    "1110101111110101",
    "1110100101010011",
    "1110100000011111",
    "1110100001001000",
    "1110100110111001",
    "1110110010101100",
    "1111000101110111",
    "1111100000010100",
    "1111111111011110",
    "1111100001001000",
    "1111000110011010",
    "1110110011100111",
    "1110101001101111",
    "1110100111010001",
    "1110101000101010",
    "1110101001101101",
    "1110100111001101",
    "1110011111110001",
    "1110010100100100",
    "1110001000010101",
    "1101111110000010",
    "1101110111110010",
    "1101110110001110",
    "1101111000101000",
    "1101111101010100",
    "1110000100110110",
    "1110010010101111",
    "1110101001111010",
    "1111001010001100",
    "1111101111101000",
    "1111101100010000",
    "1111001111100100",
    "1110111110010100",
    "1110111001000110",
    "1110111011110011",
    "1111000000011100",
    "1111000001111001",
    "1110111101000010",
    "1110110010001101",
    "1110100011110100",
    "1110010101101111",
    "1110001110110011",
    "1110010101000011",
    "1110101010011110",
    "1111001101000111",
    "1111110101010110",
    "1111100111011110",
    "1111010011000000",
    "1111010011010111",
    "1111100111010111",
    "1111111001001110",
    "1111011001001100",
    "1111000001111110",
    "1110111000010001",
    "1110111010010001",
    "1111000010011001",
    "1111001010001100",
    "1111001101001010",
    "1111001011010011",
    "1111000111110101",
    "1111000110011000",
    "1111001001010000",
    "1111010000010001",
    "1111011000110000",
    "1111100001100001",
    "1111101011110001",
    "1111111001001110",
    "1111110101010110",
    "1111100001011100",
    "1111001110100100",
    "1111000000011001",
    "1110111010100000",
    "1110111111111011",
    "1111010000110011",
    "1111101001110100",
    "1111111011101101",
    "1111100110111111",
    "1111011011100001",
    "1111011000110111",
    "1111011011111010",
    "1111100000000010",
    "1111100001101011",
    "1111011111111011",
    "1111011100100000",
    "1111011010011000",
    "1111011100000100",
    "1111100001011110",
    "1111101000101101",
    "1111101111101011",
    "1111110101001100",
    "1111111000110100",
    "1111111010010100",
    "1111111001100011",
    "1111110110111101",
    "1111110011011001",
    "1111101111101100",
    "1111101100100011",
    "1111101001110000",
    "1111101000011101",
    "1111101100111110",
    "1111111010110100",
    "1111101101110110",
    "1111010000010100",
    "1110110010110001",
    "1110011011000110",
    "1110001110001001",
    "1110010000011010",
    "1110100010111001",
    "1111000001110001",
    "1111100101001110",
    "1111111101101000",
    "1111101111101000",
    "1111110100000001",
    "1111110111001110",
    "1111011010001001",
    "1110111111010010",
    "1110101110101011",
    "1110101011100101",
    "1110110011010000",
    "1110111111010010",
    "1111001001101101",
    "1111010000001101",
    "1111010101101110",
    "1111011111001100",
    "1111110000001011",
    "1111110110011101",
    "1111011000011101",
    "1110111100010111",
    "1110101001011011",
    "1110100100001101",
    "1110101011010110",
    "1110111001000100",
    "1111000110111110",
    "1111010000011100",
    "1111010100100100",
    "1111010100011000",
    "1111010010011100",
    "1111010100101100",
    "1111100000111001",
    "1111111000111111",
    "1111100101000001",
    "1110111111001100",
    "1110011100111111",
    "1110000100111100",
    "1101111011010100",
    "1101111111110011",
    "1110001110000100",
    "1110100000011110",
    "1110110001101011",
    "1110111101110000",
    "1111000100011010",
    "1111001001101111",
    "1111010011100111",
    "1111100110010000",
    "1111111110010101",
    "1111011111000101",
    "1111000011001010",
    "1110110001001010",
    "1110101100101010",
    "1110110011001000",
    "1110111101100001",
    "1111000110000110",
    "1111001100101000",
    "1111010101000011",
    "1111100011110001",
    "1111111010101011",
    "1111100111111110",
    "1111001001011000",
    "1110110000111001",
    "1110100101101001",
    "1110101001110000",
    "1110111010010110",
    "1111010011101001",
    "1111110010000101",
    "1111101101100111",
    "1111001101111011",
    "1110110010001011",
    "1110011101111111",
    "1110010100001011",
    "1110010111010000",
    "1110100110000100",
    "1110111011100110",
    "1111010001111110",
    "1111100011111000",
    "1111101110001100",
    "1111110001011011",
    "1111101111101011",
    "1111101100000001",
    "1111101011100111",
    "1111110010110111",
    "1111111100011001",
    "1111100011001000",
    "1111000110000000",
    "1110101011110101",
    "1110011010011000",
    "1110010101111011",
    "1110011111011111",
    "1110110011110001",
    "1111001101010100",
    "1111100110000000",
    "1111111000010000",
    "1111111101011000",
    "1111110111010100",
    "1111101111011011",
    "1111100000101011",
    "1111001010001100",
    "1110101111111011",
    "1110011000000001",
    "1110001001000110",
    "1110000111101100",
    "1110010010111001",
    "1110100101001011",
    "1110110111111100",
    "1111000101101110",
    "1111001100001001",
    "1111001100000001",
    "1111000111111111",
    "1111000110011000",
    "1111001110011110",
    "1111100011010111",
    "1111111100011010",
    "1111010111000100",
    "1110110101010101",
    "1110011110001100",
    "1110010101011101",
    "1110011010101000",
    "1110101000100010",
    "1110111000101000",
    "1111000110110110",
    "1111010011011000",
    "1111100001010100",
    "1111110011011101",
    "1111110110000000",
    "1111011101100001",
    "1111000111100000",
    "1110111001001011",
    "1110110101101111",
    "1110111100010001",
    "1111001000100010",
    "1111010101001001",
    "1111011101100000",
    "1111100000001100",
    "1111011110101110",
    "1111011011011000",
    "1111011000010001",
    "1111010110010011",
    "1111010100111011",
    "1111010011001101",
    "1111010010010101",
    "1111010101011000",
    "1111011110110110",
    "1111101111011111",
    "1111111011001011",
    "1111100110110001",
    "1111011000101010",
    "1111010100010010",
    "1111011001011000",
    "1111100011010000",
    "1111101100000010",
    "1111101110111011",
    "1111101001100011",
    "1111011101001110",
    "1111001100100110",
    "1110111011110101",
    "1110110010001000",
    "1110110101100000",
    "1111000111101010",
    "1111100110010011",
    "1111110101100000",
    "1111010100010111",
    "1110111101010001",
    "1110110100101111",
    "1110111010001110",
    "1111001000101000",
    "1111011001010101",
    "1111100101111100",
    "1111101010100100",
    "1111100111001010",
    "1111011101110111",
    "1111010001111110",
    "1111001000001110",
    "1111000101110110",
    "1111001110010111",
    "1111100001110110",
    "1111111100101001",
    "1111100111011100",
    "1111010000011111",
    "1111000010100111",
    "1110111111100011",
    "1111000100101110",
    "1111001100011001",
    "1111010001001101",
    "1111010000000101",
    "1111001001110101",
    "1111000001110110",
    "1110111010111100",
    "1110111000010110",
    "1110111110000101",
    "1111001101111000",
    "1111100110100100",
    "1111111011110110",
    "1111011111110110",
    "1111001010110100",
    "1110111111100110",
    "1110111110101110",
    "1111000100101010",
    "1111001100000100",
    "1111010000100100",
    "1111001111101001",
    "1111001100010100",
    "1111001110001001",
    "1111011011000010",
    "1111110101011011",
    "1111100101100111",
    "1110111110011011",
    "1110011101011011",
    "1110001001100101",
    "1110001000010110",
    "1110011010100000",
    "1110111011110010",
    "1111100101000001",
    "1111110010000000",
    "1111010000011100",
    "1110111010111100",
    "1110110100011000",
    "1110111011011000",
    "1111001010001100",
    "1111011010100110",
    "1111100111010010",
    "1111101110010101",
    "1111110010110011",
    "1111111001001110",
    "1111111010101001",
    "1111100111000101",
    "1111001110001101",
    "1110110101100111",
    "1110100011111011",
    "1110011110101110",
    "1110100111010000",
    "1110111001101101",
    "1111010000010010",
    "1111100110111001",
    "1111111101101000",
    "1111101001010111",
    "1111001100111101",
    "1110101110000101",
    "1110010000011010",
    "1101111001111001",
    "1101110000100011",
    "1101110111011111",
    "1110001100100110",
    "1110101001110101",
    "1111000111101101",
    "1111011111100110",
    "1111101111111101",
    "1111111100101101",
    "1111110100100001",
    "1111011111101011",
    "1111000100100111",
    "1110101001010011",
    "1110010110101100",
    "1110010100101100",
    "1110100110101000",
    "1111001000110100",
    "1111110010111000",
    "1111100100011111",
    "1111000101010010",
    "1110110011100010",
    "1110110000111000",
    "1110111101000010",
    "1111010101010011",
    "1111110101010110",
    "1111101000000101",
    "1111001001011001",
    "1110110100011101",
    "1110101101001111",
    "1110110101000011",
    "1111001000111100",
    "1111100010110110",
    "1111111100011100",
    "1111101110101010",
    "1111011111001000",
    "1111010011010011",
    "1111001001011000",
    "1110111111111101",
    "1110110111010110",
    "1110110001100010",
    "1110110000011001",
    "1110110100011000",
    "1110111100010110",
    "1111000101111011",
    "1111001110101110",
    "1111010110100000",
    "1111100000110110",
    "1111110010110101",
    "1111110001010010",
    "1111001101011011",
    "1110100111111110",
    "1110001001011110",
    "1101111001000110",
    "1101111010100101",
    "1110001011010001",
    "1110100011011010",
    "1110111010000111",
    "1111001001001110",
    "1111010001110100",
    "1111011010010100",
    "1111101000001110",
    "1111111101111110",
    "1111100110111100",
    "1111001101011110",
    "1110111100110010",
    "1110111010001001",
    "1111000101001001",
    "1111011000011010",
    "1111101111011001",
    "1111111000111110",
    "1111100010010101",
    "1111001100101101",
    "1110111001111010",
    "1110101100011001",
    "1110100110001110",
    "1110101001001011",
    "1110110100001000",
    "1111000010110011",
    "1111010001100001",
    "1111100000000111",
    "1111110001100011",
    "1111110111011000",
    "1111011010101011",
    "1110111011100110",
    "1110100000011001",
    "1110010000100111",
    "1110010001111110",
    "1110100100101100",
    "1111000011001010",
    "1111100101000000",
    "1111111011110100",
    "1111100000011111",
    "1111000110100111",
    "1110101011111100",
    "1110010000101001",
    "1101111000010101",
    "1101101000011000",
    "1101100101100101",
    "1101110001001100",
    "1110000110110001",
    "1110100000110110",
    "1110111100101011",
    "1111011000111100",
    "1111110101111010",
    "1111101100100001",
    "1111010001000000",
    "1110111010011011",
    "1110101100100011",
    "1110101010010110",
    "1110110010010000",
    "1111000000000111",
    "1111001110101110",
    "1111011001001100",
    "1111011101011001",
    "1111011100101110",
    "1111011100101101",
    "1111100100110111",
    "1111111000110110",
    "1111101001011001",
    "1111001000011000",
    "1110101100110000",
    "1110011101101000",
    "1110011110000101",
    "1110101011111101",
    "1111000000110001",
    "1111010101011111",
    "1111100100110011",
    "1111101100010110",
    "1111101100110000",
    "1111101001101101",
    "1111101001011111",
    "1111110001001100",
    "1111111101101110",
    "1111100110010000",
    "1111001110010111",
    "1110111100000100",
    "1110110011101110",
    "1110110110001001",
    "1111000000000011",
    "1111001100100001",
    "1111010110110110",
    "1111011011100000",
    "1111011001110100",
    "1111010010111110",
    "1111001001101011",
    "1111000001100001",
    "1110111100101011",
    "1110111011010110",
    "1110111100100011",
    "1110111110101101",
    "1111000000001111",
    "1111000001001100",
    "1111000100111110",
    "1111010000000010",
    "1111100100001101",
    "1111111111110111",
    "1111100000110011",
    "1111000100011111",
    "1110110000001111",
    "1110101000000110",
    "1110101011111010",
    "1110110111000011",
    "1111000011101100",
    "1111001100101101",
    "1111001111100001",
    "1111001110010110",
    "1111001111001101",
    "1111011000100000",
    "1111101101100000",
    "1111110011111100",
    "1111010010110100",
    "1110110111000110",
    "1110100111001110",
    "1110100110000100",
    "1110110000100110",
    "1110111111111011",
    "1111001101011110",
    "1111010100111100",
    "1111010101101100",
    "1111010001110100",
    "1111001100010110",
    "1111001000011101",
    "1111001000000110",
    "1111001101001010",
    "1111011001111010",
    "1111101110100111",
    "1111110110010101",
    "1111011001011000",
    "1111000011000101",
    "1110111100001001",
    "1111001001101011",
    "1111101010010011",
    "1111101011011000",
    "1111000011111110",
    "1110101010001001",
    "1110100011111100",
    "1110101111010001",
    "1111000100001000",
    "1111011001011110",
    "1111101010000101",
    "1111110111100010",
    "1111111001000111",
    "1111100100011010",
    "1111001010010011",
    "1110101111001111",
    "1110011010000111",
    "1110010001011010",
    "1110010111101000",
    "1110101001101000",
    "1111000000010100",
    "1111010101010101",
    "1111100111110101",
    "1111111011110010",
    "1111101010100000",
    "1111001010001011",
    "1110100111011010",
    "1110001001110111",
    "1101111001100000",
    "1101111011010100",
    "1110001110001001",
    "1110101011000001",
    "1111001001001001",
    "1111100010101110",
    "1111111000111001",
    "1111101111000010",
    "1111010000111000",
    "1110101011111111",
    "1110000101000001",
    "1101100100000110",
    "1101010001001000",
    "1101010000101001",
    "1101100000110110",
    "1101111010110100",
    "1110010110001110",
    "1110101100001111",
    "1110111010011001",
    "1111000010010010",
    "1111000110011101",
    "1111001001001011",
    "1111001011010011",
    "1111001100010100",
    "1111001011100110",
    "1111001000111110",
    "1111000101000110",
    "1111000001011110",
    "1110111111100001",
    "1110111111100011",
    "1111000000001010",
    "1110111111001010",
    "1110111011011101",
    "1110111000001110",
    "1110111011111100",
    "1111001011101010",
    "1111101000110110",
    "1111110000010101",
    "1111000111111001",
    "1110100110010110",
    "1110010010110001",
    "1110001111001100",
    "1110010111001011",
    "1110100011111000",
    "1110101111010001",
    "1110110110001000",
    "1110111001010001",
    "1110111011001100",
    "1110111101110101",
    "1111000011100010",
    "1111001110110101",
    "1111100000011111",
    "1111110111010100",
    "1111101111101110",
    "1111011001000010",
    "1111001000010000",
    "1111000000000000",
    "1111000001101110",
    "1111001100110000",
    "1111100000001111",
    "1111111010111000",
    "1111100101111100",
    "1111000101101010",
    "1110101000101100",
    "1110010011111100",
    "1110001010010001",
    "1110001100110010",
    "1110011001100010",
    "1110101011110000",
    "1111000001000010",
    "1111011000111111",
    "1111110011000010",
    "1111110001101100",
    "1111011000100111",
    "1111000101100101",
    "1110111011100000",
    "1110111100111000",
    "1111001001000110",
    "1111011010110100",
    "1111101100110011",
    "1111111101011011",
    "1111110001011101",
    "1111011100101110",
    "1111000010111101",
    "1110100110001110",
    "1110001011010100",
    "1101111000011110",
    "1101110011001000",
    "1101111011111111",
    "1110001111000000",
    "1110100101111110",
    "1110111010011001",
    "1111001010100101",
    "1111011010011000",
    "1111101110000111",
    "1111110111111100",
    "1111011001100000",
    "1110111100111101",
    "1110101010001110",
    "1110101001000111",
    "1110111110010001",
    "1111100110001101",
    "1111101000110110",
    "1110111010110010",
    "1110011001010001",
    "1110001000100000",
    "1110001000010110",
    "1110010101101100",
    "1110101010010110",
    "1110111111011100",
    "1111001111110110",
    "1111011001000110",
    "1111011011100001",
    "1111011001011101",
    "1111010101011010",
    "1111010011111000",
    "1111011011100110",
    "1111110001001000",
    "1111101011111000",
    "1111000001011001",
    "1110011001001011",
    "1101111100100110",
    "1101110010011100",
    "1101111100100011",
    "1110010111001001",
    "1110111101010110",
    "1111101010000101",
    "1111100111111111",
    "1110111101001010",
    "1110011001101111",
    "1110000010100001",
    "1101111010110010",
    "1110000100011000",
    "1110011111010001",
    "1111001000010000",
    "1111111001100010",
    "1111010100001011",
    "1110101001001001",
    "1110001011111100",
    "1101111111110001",
    "1110000011010111",
    "1110010001100110",
    "1110100011101111",
    "1110110100101111",
    "1111000100001010",
    "1111010101010101",
    "1111101011100010",
    "1111111001000010",
    "1111011011111111",
    "1111000010100111",
    "1110110010011001",
    "1110101111000111",
    "1110110111110100",
    "1111000111001101",
    "1111010110111111",
    "1111100010000110",
    "1111100111001101",
    "1111101011011000",
    "1111110110011011",
    "1111110010100010",
    "1111001111110011",
    "1110101000100011",
    "1110000111010011",
    "1101110100111001",
    "1101110110011000",
    "1110001011010100",
    "1110101111100100",
    "1111011101101011",
    "1111110000101001",
    "1111000001100111",
    "1110011010101010",
    "1110000000100011",
    "1101110110000011",
    "1101111010110000",
    "1110001011100000",
    "1110100010010000",
    "1110111000100010",
    "1111001001110101",
    "1111010100010111",
    "1111011000101100",
    "1111011001001110",
    "1111011001011011",
    "1111011100100000",
    "1111100011010101",
    "1111101101000011",
    "1111111001000001",
    "1111110111111100",
    "1111100100110100",
    "1111001101011001",
    "1110110011011101",
    "1110011011100101",
    "1110001011000111",
    "1110000110001001",
    "1110001101100011",
    "1110011101100100",
    "1110101111101001",
    "1110111101000100",
    "1111000001010100",
    "1110111011110111",
    "1110101111101000",
    "1110100001000101",
    "1110010101000110",
    "1110001111001000",
    "1110001111110101",
    "1110010101101111",
    "1110011110011110",
    "1110101000010101",
    "1110110010100010",
    "1110111101101001",
    "1111001100100110",
    "1111100010000101",
    "1111111110010101",
    "1111100001000111",
    "1111000001110000",
    "1110101001101000",
    "1110011101010001",
    "1110011110101001",
    "1110101011000110",
    "1110111101001110",
    "1111010000010111",
    "1111100000110000",
    "1111101100001111",
    "1111110010101110",
    "1111110100100100",
    "1111110010111010",
    "1111101111000101",
    "1111101010000011",
    "1111100110010010",
    "1111100111010110",
    "1111101111001011",
    "1111111101010001",
    "1111110001010110",
    "1111100001010000",
    "1111010110011000",
    "1111010011011010",
    "1111011000101111",
    "1111100011111100",
    "1111110001011100",
    "1111111110101001",
    "1111110100111011",
    "1111101000011001",
    "1111011011010100",
    "1111001111000010",
    "1111000101101110",
    "1111000001000010",
    "1111000001010111",
    "1111000101100101",
    "1111001011000001",
    "1111001111110110",
    "1111010110001011",
    "1111100001111110",
    "1111110110000001",
    "1111101101110010",
    "1111001101111010",
    "1110110001000111",
    "1110011110001001",
    "1110011001110000",
    "1110100010111001",
    "1110110011101001",
    "1111000111001101",
    "1111011100000010",
    "1111110010101001",
    "1111110011110000",
    "1111011000010000",
    "1110111110010111",
    "1110101010110111",
    "1110100011100001",
    "1110101011000110",
    "1110111110110101",
    "1111011000110100",
    "1111110001111001",
    "1111111001111100",
    "1111101000101010",
    "1111010110010110",
    "1111000000011001",
    "1110100111010110",
    "1110010000100100",
    "1110000010111001",
    "1110000011010000",
    "1110010010110011",
    "1110101100100110",
    "1111001000000001",
    "1111011101010110",
    "1111101000000111",
    "1111101001001010",
    "1111100100100100",
    "1111011110011011",
    "1111011001110111",
    "1111010111111010",
    "1111010111010011",
    "1111010110010010",
    "1111010011010111",
    "1111001111011010",
    "1111001111001010",
    "1111010111000110",
    "1111100111110111",
    "1111111101100001",
    "1111101110111101",
    "1111100011100100",
    "1111100001101011",
    "1111100101110110",
    "1111101000110011",
    "1111100011101001",
    "1111010100000001",
    "1110111100110000",
    "1110100100011100",
    "1110010010011001",
    "1110001010111100",
    "1110001110000101",
    "1110011000101000",
    "1110100101110111",
    "1110110010101100",
    "1110111110101000",
    "1111001011011110",
    "1111011011101111",
    "1111110000011001",
    "1111111000101000",
    "1111100100001010",
    "1111010110111111",
    "1111010011011010",
    "1111010111100000",
    "1111011110011111",
    "1111100010111001",
    "1111100000111101",
    "1111011000010110",
    "1111001011100001",
    "1110111110010001",
    "1110110011111011",
    "1110101110001101",
    "1110101100110010",
    "1110101101101101",
    "1110110000000011",
    "1110110110101010",
    "1111000101010000",
    "1111011101110011",
    "1111111111000001",
    "1111011100101101",
    "1110111101000101",
    "1110101000110100",
    "1110100011001011",
    "1110101001100011",
    "1110110100111011",
    "1110111110001010",
    "1111000000100100",
    "1110111011100000",
    "1110110010000101",
    "1110101001111101",
    "1110101001101111",
    "1110110101010000",
    "1111001011111101",
    "1111101001101111",
    "1111110111011000",
    "1111011101001111",
    "1111001011100110",
    "1111000011101001",
    "1111000011100100",
    "1111001000011110",
    "1111001111111000",
    "1111010111100000",
    "1111011110011001",
    "1111100110001101",
    "1111110001010001",
    "1111111111100001",
    "1111101110011010",
    "1111100000101100",
    "1111011100001110",
    "1111100101000011",
    "1111111011111010",
    "1111100011111000",
    "1111000011001011",
    "1110101100001110",
    "1110101000001000",
    "1110111010101101",
    "1111100001001101",
    "1111101100011111",
    "1110111010100101",
    "1110010100100101",
    "1110000001010000",
    "1110000001100110",
    "1110010000001101",
    "1110100100011100",
    "1110110110011000",
    "1111000001011111",
    "1111000111110010",
    "1111001111011001",
    "1111011101000100",
    "1111110010111010",
    "1111110001010111",
    "1111010101101110",
    "1111000000000111",
    "1110110101010111",
    "1110110101101111",
    "1110111101101000",
    "1111001010111111",
    "1111011101010100",
    "1111110100100001",
    "1111101111110011",
    "1111010011011010",
    "1110111011011011",
    "1110101100010011",
    "1110101010000010",
    "1110110100011000",
    "1111000110110010",
    "1111011110101011",
    "1111111011000001",
    "1111100101000001",
    "1111000010110110",
    "1110100010011101",
    "1110001000110101",
    "1101111010011110",
    "1101111011010011",
    "1110001100001001",
    "1110101011011001",
    "1111010110001110",
    "1111111000110000",
    "1111001000010011",
    "1110011110100110",
    "1110000000100100",
    "1101110000011010",
    "1101101101111000",
    "1101110110111011",
    "1110000111010001",
    "1110011001111010",
    "1110101010101101",
    "1110110111001011",
    "1110111110110000",
    "1111000010001000",
    "1111000011001011",
    "1111000100001011",
    "1111000111101100",
    "1111010001101011",
    "1111100101000001",
    "1111111111000000",
    "1111011110110101",
    "1111000001110100",
    "1110101111010010",
    "1110101100010001",
    "1110111001100010",
    "1111010001110000",
    "1111101011111001",
    "1111111111111110",
    "1111110110111011",
    "1111111001000101",
    "1111111111011000",
    "1111111010011110",
    "1111111101110001",
    "1111110101010111",
    "1111100011001000",
    "1111010010001000",
    "1111001000010000",
    "1111001001000111",
    "1111010011010101",
    "1111100000100111",
    "1111101010011101",
    "1111101101010000",
    "1111101001000100",
    "1111100001100110",
    "1111011011010100",
    "1111011001110111",
    "1111011110110101",
    "1111101000000111",
    "1111110001110010",
    "1111111000011100",
    "1111111001101010",
    "1111110101110011",
    "1111110001011111",
    "1111110011010001",
    "1111111111010111",
    "1111101010001000",
    "1111001101101110",
    "1110110010010000",
    "1110011101111010",
    "1110010101010000",
    "1110011001000100",
    "1110100110000000",
    "1110110111000110",
    "1111000111000011",
    "1111010001111011",
    "1111010110110001",
    "1111010110000000",
    "1111010010101111",
    "1111010011011100",
    "1111011101000111",
    "1111110001001000",
    "1111110011001111",
    "1111010110101101",
    "1111000000001101",
    "1110110100111011",
    "1110110111010001",
    "1111000100010000",
    "1111010101011101",
    "1111100100100100",
    "1111101100110000",
    "1111101101010110",
    "1111101011011010",
    "1111101110101011",
    "1111111101010100",
    "1111100111001101",
    "1111000100000000",
    "1110100001100111",
    "1110001000001110",
    "1101111110001001",
    "1110000011110110",
    "1110010011110001",
    "1110101001000100",
    "1111000001111000",
    "1111011101100000",
    "1111111011101100",
    "1111100110001101",
    "1111001100011011",
    "1110111010010100",
    "1110110011010000",
    "1110110111111111",
    "1111000100011111",
    "1111010011010011",
    "1111100001010000",
    "1111101110111111",
    "1111111111001100",
    "1111101100001111",
    "1111010100011000",
    "1110111101001010",
    "1110101100101010",
    "1110101000011010",
    "1110110010000010",
    "1111000101110010",
    "1111011100101000",
    "1111101111001100",
    "1111111011001111",
    "1111111011011101",
    "1111110000010101",
    "1111100001000011",
    "1111001111100100",
    "1111000001110011",
    "1110111101101101",
    "1111000110101111",
    "1111011011111100",
    "1111110111011001",
    "1111101110010101",
    "1111011010010011",
    "1111001011101010",
    "1110111101001100",
    "1110101010100101",
    "1110010011001000",
    "1101111010001100",
    "1101100110000110",
    "1101011101100000",
    "1101100100011000",
    "1101111001011001",
    "1110010110010110",
    "1110110011111000",
    "1111001101011110",
    "1111100011011101",
    "1111111001001000",
    "1111101111001000",
    "1111010101001000",
    "1110111010100010",
    "1110100010110001",
    "1110010001101001",
    "1110001001001100",
    "1110001000111111",
    "1110001110100001",
    "1110010110110100",
    "1110011111101110",
    "1110101000100101",
    "1110110001100110",
    "1110111010011101",
    "1111000010011100",
    "1111001000100111",
    "1111001100010110",
    "1111001111001100",
    "1111010100111011",
    "1111100000111110",
    "1111110100000111",
    "1111110011111100",
    "1111011011110101",
    "1111001000000110",
    "1110111011101101",
    "1110110110110001",
    "1110110110010011",
    "1110110110100010",
    "1110110101001110",
    "1110110010010000",
    "1110101110111011",
    "1110101100110011",
    "1110101100110010",
    "1110101111010010",
    "1110110011101010",
    "1110111000010101",
    "1110111100000100",
    "1110111110111000",
    "1111000001001010",
    "1111000100111001",
    "1111001110100100",
    "1111100001101110",
    "1111111110101001",
    "1111011110001100",
    "1110111011101011",
    "1110100000101011",
    "1110010010001011",
    "1110010010010000",
    "1110011101110111",
    "1110101110001101",
    "1110111100011011",
    "1111000011101111",
    "1111000011010010",
    "1110111111101000",
    "1111000000011111",
    "1111001100100000",
    "1111100101111100",
    "1111110110111001",
    "1111010001110000",
    "1110110010100110",
    "1110011111110011",
    "1110011011100101",
    "1110100010011001",
    "1110101110000000",
    "1110111000101101",
    "1110111111100011",
    "1111000011011000",
    "1111000110101010",
    "1111001010111000",
    "1111010000011111",
    "1111010101100111",
    "1111010110111111",
    "1111010010100111",
    "1111001000011011",
    "1110111011011101",
    "1110110000011110",
    "1110101011101000",
    "1110110001011010",
    "1111000101001000",
    "1111100110010000",
    "1111101110110100",
    "1111000000111000",
    "1110010111110101",
    "1101111010000010",
    "1101101011100000",
    "1101101100001111",
    "1101110111010011",
    "1110000110001001",
    "1110010011000001",
    "1110011010100101",
    "1110011100100110",
    "1110011010111000",
    "1110011000011010",
    "1110011000010101",
    "1110011100010001",
    "1110100100010010",
    "1110101111011111",
    "1110111110010111",
    "1111010011001000",
    "1111101111010110",
    "1111101101110000",
    "1111001000101010",
    "1110101000100010",
    "1110010100010111",
    "1110010000011010",
    "1110011100011100",
    "1110110010111110",
    "1111001100000111",
    "1111100010101111",
    "1111110110101000",
    "1111110101111011",
    "1111100001000010",
    "1111001011001110",
    "1110110111010000",
    "1110101000101111",
    "1110100011010111",
    "1110100111111010",
    "1110110010111110",
    "1110111111001111",
    "1111000111010000",
    "1111001001001011",
    "1111001010000100",
    "1111010000110000",
    "1111100001100010",
    "1111111100000011",
    "1111100111000110",
    "1111010010101001",
    "1111001111010100",
    "1111100001001100",
    "1111111100010000",
    "1111010100000110",
    "1110110001111110",
    "1110100000100001",
    "1110100101001011",
    "1110111110010001",
    "1111100110000001",
    "1111101100100010",
    "1111000010111000",
    "1110100010111000",
    "1110010000001100",
    "1110001011010001",
    "1110010000100100",
    "1110011011111101",
    "1110101001101111",
    "1110110110010101",
    "1110111111110000",
    "1111000101000001",
    "1111000110101101",
    "1111001001001100",
    "1111010010110100",
    "1111100111110101",
    "1111110111000101",
    "1111001110101001",
    "1110100111010001",
    "1110001000101000",
    "1101111000000110",
    "1101110110111001",
    "1110000000110001",
    "1110001111011010",
    "1110011101011100",
    "1110100111101111",
    "1110101110110101",
    "1110110101000001",
    "1110111100010110",
    "1111000101111001",
    "1111010001101100",
    "1111100000011010",
    "1111110011011101",
    "1111110101000000",
    "1111011010011000",
    "1111000000011111",
    "1110101101111000",
    "1110101001110100",
    "1110111000111100",
    "1111011001110101",
    "1111111011100110",
    "1111010010001011",
    "1110110011111000",
    "1110100110011000",
    "1110101001101011",
    "1110111010110010",
    "1111010101111110",
    "1111110110101011",
    "1111100111001111",
    "1111000111110010",
    "1110101110111010",
    "1110011111001010",
    "1110011010000100",
    "1110011111101100",
    "1110101101001010",
    "1110111101110101",
    "1111001101101000",
    "1111011001100011",
    "1111100001011010",
    "1111101000100011",
    "1111110011011011",
    "1111111010110110",
    "1111100011000001",
    "1111001010010100",
    "1110110111001000",
    "1110101110100110",
    "1110110011000101",
    "1111000010000011",
    "1111010101010011",
    "1111100111000100",
    "1111110011110101",
    "1111111011001111",
    "1111111111011011",
    "1111111100111010",
    "1111110111011110",
    "1111101111110001",
    "1111100111110110",
    "1111100001010100",
    "1111011100010011",
    "1111011000001011",
    "1111010011101100",
    "1111001101111111",
    "1111000111101111",
    "1111000011000001",
    "1111000010101110",
    "1111001000010101",
    "1111010010100001",
    "1111011110010111",
    "1111101000101110",
    "1111101111001000",
    "1111110001001101",
    "1111110010001000",
    "1111110111100101",
    "1111111010001000",
    "1111100010111101",
    "1111000111001001",
    "1110101110011100",
    "1110100000010101",
    "1110100010000110",
    "1110110110011011",
    "1111011011000010",
    "1111110110101010",
    "1111000111001001",
    "1110011111000100",
    "1110000100011010",
    "1101111001010011",
    "1101111101101101",
    "1110010000011010",
    "1110101110010110",
    "1111010010111101",
    "1111111000010101",
    "1111100111110101",
    "1111010010100010",
    "1111001010010100",
    "1111001111010010",
    "1111011111010100",
    "1111110110111101",
    "1111101101101110",
    "1111010010110001",
    "1110111011000100",
    "1110101000110010",
    "1110011110001100",
    "1110011100111000",
    "1110100100000000",
    "1110110000001000",
    "1110111101100011",
    "1111001011000111",
    "1111011010110101",
    "1111101110111000",
    "1111111000111001",
    "1111011111001100",
    "1111000111101100",
    "1110110101101111",
    "1110101011110010",
    "1110101001111101",
    "1110101101101011",
    "1110110011010011",
    "1110111000010110",
    "1110111100001100",
    "1110111111101110",
    "1111000100000011",
    "1111001001010110",
    "1111001111011111",
    "1111010110110100",
    "1111100000111011",
    "1111101111111011",
    "1111111011101011",
    "1111100011111000",
    "1111001101001110",
    "1110111101110111",
    "1110111011011011",
    "1111001000101000",
    "1111100010110001",
    "1111111101011010",
    "1111100000001111",
    "1111001011111000",
    "1111000010111011",
    "1111000100010011",
    "1111001100010111",
    "1111010101101010",
    "1111011011011110",
    "1111011011111100",
    "1111010111111100",
    "1111010001111101",
    "1111001100010001",
    "1111001000000110",
    "1111000101011111",
    "1111000011101111",
    "1111000010000010",
    "1110111111110001",
    "1110111101011100",
    "1110111101010001",
    "1111000010011010",
    "1111001110101000",
    "1111100001001010",
    "1111110111011000",
    "1111110001111111",
    "1111011101111010",
    "1111001110001010",
    "1111000011000101",
    "1110111011100001",
    "1110110101110100",
    "1110110001000000",
    "1110101111001100",
    "1110110100011101",
    "1111000011100001",
    "1111011011110111",
    "1111111001110101",
    "1111101000011010",
    "1111010000111000",
    "1111000100010000",
    "1111000011110110",
    "1111001100011100",
    "1111011001101011",
    "1111101010000001",
    "1111111110100000",
    "1111100111001111",
    "1111000111110111",
    "1110100111011011",
    "1110001011100101",
    "1101111010001110",
    "1101111000000100",
    "1110000100101010",
    "1110011011100110",
    "1110111001011000",
    "1111011011101000",
    "1111111111010000",
    "1111011000110111",
    "1110110100110110",
    "1110011000001100",
    "1110000111101010",
    "1110000111011101",
    "1110010111011010",
    "1110110001110110",
    "1111001111011110",
    "1111101000011001",
    "1111111000001110",
    "1111111110001000",
    "1111110100011100",
    "1111100100110100",
    "1111001101010001",
    "1110110100011000",
    "1110100100110110",
    "1110100111100000",
    "1111000000010101",
    "1111101001110110",
    "1111101000011001",
    "1111000011100010",
    "1110110000111011",
    "1110110010000110",
    "1111000011100110",
    "1111100000100111",
    "1111111101001001",
    "1111011011010001",
    "1110111101001111",
    "1110100110001101",
    "1110010111100011",
    "1110010001111000",
    "1110010100110111",
    "1110011101101000",
    "1110101010000100",
    "1110111010110111",
    "1111010000101011",
    "1111101011100001",
    "1111110110011000",
    "1111011001010011",
    "1111000001001100",
    "1110110010001101",
    "1110101111100100",
    "1110110111110001",
    "1111000110000001",
    "1111010101000101",
    "1111100000000101",
    "1111100111000011",
    "1111101111100001",
    "1111111111010000",
    "1111100110010010",
    "1111000011010010",
    "1110011111110101",
    "1110000100101010",
    "1101111000111010",
    "1101111111101100",
    "1110010101010000",
    "1110110001111011",
    "1111001101111000",
    "1111100010110100",
    "1111101111111100",
    "1111111010000100",
    "1111111001000011",
    "1111100101110100",
    "1111001101000100",
    "1110110101001000",
    "1110100101011000",
    "1110100011010011",
    "1110110001101100",
    "1111001111011110",
    "1111110111011000",
    "1111011101010110",
    "1110110101101110",
    "1110010111101100",
    "1110000110111001",
    "1110000101010010",
    "1110010001111110",
    "1110101000010000",
    "1111000001100111",
    "1111011001011001",
    "1111101111101011",
    "1111111000001000",
    "1111011011011110",
    "1110111010111101",
    "1110011010110000",
    "1110000000100111",
    "1101110010100110",
    "1101110101000000",
    "1110000111000100",
    "1110100011010010",
    "1111000001111011",
    "1111011011110111",
    "1111101100110110",
    "1111110100110001",
    "1111110110000001",
    "1111110100011001",
    "1111110010110110",
    "1111110001111001",
    "1111110000110101",
    "1111110000000001",
    "1111110001110001",
    "1111111000110001",
    "1111111001100010",
    "1111100110011000",
    "1111010001110001",
    "1111000000101110",
    "1110110111100111",
    "1110111001011000",
    "1111000111000001",
    "1111011111010010",
    "1111111101111110",
    "1111100010100110",
    "1111000111101100",
    "1110110101001101",
    "1110101100111100",
    "1110101110000111",
    "1110110101110110",
    "1111000000001101",
    "1111001001100111",
    "1111001111110000",
    "1111010010010000",
    "1111010010001011",
    "1111010010110001",
    "1111011000111110",
    "1111101000100011",
    "1111111110111101",
    "1111100010110110",
    "1111001011001010",
    "1110111111001000",
    "1111000010010111",
    "1111010011100001",
    "1111101100100000",
    "1111111001111111",
    "1111100110000110",
    "1111011100001001",
    "1111011110001111",
    "1111101100001000",
    "1111111100100101",
    "1111100000011010",
    "1111000100001000",
    "1110101011110011",
    "1110011010101011",
    "1110010010011100",
    "1110010010100010",
    "1110011000110100",
    "1110100010010101",
    "1110101100001010",
    "1110110101001101",
    "1111000000011001",
    "1111010001111011",
    "1111101100010001",
    "1111110001110010",
    "1111001110100001",
    "1110110001100111",
    "1110100001000111",
    "1110011111011010",
    "1110101001010000",
    "1110110111011011",
    "1111000011000101",
    "1111001001101010",
    "1111001110110001",
    "1111011000010110",
    "1111101010010000",
    "1111111011010000",
    "1111011100011001",
    "1110111111111000",
    "1110101100011110",
    "1110100101101001",
    "1110101010111101",
    "1110111011001110",
    "1111010100011000",
    "1111110011011101",
    "1111101010010011",
    "1111001001010001",
    "1110101110110011",
    "1110011111101000",
    "1110011111011111",
    "1110101101101001",
    "1111000101110001",
    "1111100100101010",
    "1111111000011100",
    "1111010100001010",
    "1110110001001010",
    "1110010011110110",
    "1101111111101000",
    "1101110110110110",
    "1101111011101101",
    "1110001101000000",
    "1110100101111001",
    "1111000001100100",
    "1111011101111010",
    "1111111011011100",
    "1111100100100111",
    "1111000010011111",
    "1110100000011110",
    "1110000010101001",
    "1101101110011100",
    "1101101000011101",
    "1101110001001101",
    "1110000101010101",
    "1110011111000111",
    "1110111000001000",
    "1111001100100101",
    "1111011101000100",
    "1111101101000000",
    "1111111111110010",
    "1111101001111101",
    "1111010011000011",
    "1110111111110011",
    "1110110101000101",
    "1110110110111001",
    "1111000110101000",
    "1111100001101001",
    "1111111110001101",
    "1111011111101001",
    "1111000111101010",
    "1110111001001011",
    "1110110101011011",
    "1110111011111111",
    "1111001010011110",
    "1111011101110010",
    "1111110011011101",
    "1111110110100000",
    "1111100010010000",
    "1111010010010101",
    "1111001001111101",
    "1111001011100101",
    "1111010111010011",
    "1111101010110001",
    "1111111110001111",
    "1111101000001100",
    "1111010101100111",
    "1111000111001110",
    "1110111100010111",
    "1110110011111000",
    "1110101100111101",
    "1110100111101111",
    "1110100101010011",
    "1110100110110100",
    "1110101100010001",
    "1110110100100111",
    "1111000000000101",
    "1111010000010100",
    "1111100110011111",
    "1111111101011011",
    "1111011101101001",
    "1110111110000101",
    "1110100011011101",
    "1110010010101001",
    "1110001110010100",
    "1110010100111001",
    "1110100010001010",
    "1110110000110110",
    "1110111101001001",
    "1111000111001110",
    "1111010010000000",
    "1111100000010100",
    "1111110011101101",
    "1111110101010101",
    "1111011111010100",
    "1111001111000000",
    "1111001000000110",
    "1111001010110000",
    "1111010011001111",
    "1111011100000100",
    "1111100000110000",
    "1111011111001100",
    "1111011000011011",
    "1111001111010010",
    "1111000110100100",
    "1111000001111000",
    "1111000101101111",
    "1111010100010111",
    "1111101100110001",
    "1111110101000110",
    "1111010111110001",
    "1111000001001100",
    "1110110101101111",
    "1110110111100111",
    "1111000110110100",
    "1111100001011100",
    "1111111100101011",
    "1111011001011101",
    "1110111011000001",
    "1110100110110110",
    "1110100000011001",
    "1110101000000011",
    "1110111010110111",
    "1111010010011111",
    "1111101000000110",
    "1111111001001111",
    "1111110111111000",
    "1111100111110111",
    "1111010100110011",
    "1110111111110000",
    "1110101011101101",
    "1110011100101011",
    "1110010111000110",
    "1110011100010100",
    "1110101001011110",
    "1110111001110101",
    "1111001000010110",
    "1111010011111110",
    "1111100001100010",
    "1111110110010001",
    "1111101011101100",
    "1111000110110010",
    "1110100010100111",
    "1110000111101100",
    "1101111100101101",
    "1110000100010101",
    "1110011010011000",
    "1110110110110010",
    "1111010001111000",
    "1111100110011001",
    "1111110011110010",
    "1111111100000110",
    "1111111110110010",
    "1111111011011001",
    "1111111001100011",
    "1111111010101100",
    "1111111111110011",
    "1111110110010010",
    "1111101100110001",
    "1111101010000001",
    "1111110011001100",
    "1111110111000110",
    "1111011001111101",
    "1110111101011001",
    "1110101000100011",
    "1110011111110011",
    "1110100011001000",
    "1110101110000101",
    "1110111010100101",
    "1111000101010101",
    "1111001111111010",
    "1111011101110101",
    "1111110001001001",
    "1111110111000101",
    "1111011111001100",
    "1111001100011001",
    "1111000010111011",
    "1111000100000000",
    "1111001100010110",
    "1111010110011011",
    "1111011101011011",
    "1111011111001010",
    "1111011111010001",
    "1111100100011100",
    "1111110011000001",
    "1111110100010110",
    "1111010101100100",
    "1110110111001000",
    "1110011111010110",
    "1110010010110011",
    "1110010010001111",
    "1110011010100011",
    "1110100111010001",
    "1110110100010011",
    "1110111111100110",
    "1111001001000001",
    "1111010000110101",
    "1111011000100011",
    "1111100010111101",
    "1111110001001101",
    "1111111101011101",
    "1111101011101100",
    "1111011101001001",
    "1111010101000001",
    "1111010101001001",
    "1111011101101011",
    "1111101100000011",
    "1111111011110111",
    "1111110111011100",
    "1111110000010110",
    "1111101101110101",
    "1111101100100110",
    "1111101000111110",
    "1111100000100111",
    "1111010100000101",
    "1111000110110001",
    "1110111101001010",
    "1110111010101111",
    "1111000000010010",
    "1111001011011001",
    "1111010111111100",
    "1111100100011100",
    "1111110010100100",
    "1111111011100011",
    "1111100101010101",
    "1111001101011011",
    "1110111000101101",
    "1110101011111000",
    "1110101010110000",
    "1110110101100101",
    "1111001000011010",
    "1111011110011100",
    "1111110100010000",
    "1111110111011011",
    "1111100100010000",
    "1111010010011111",
    "1111000011010101",
    "1110111000001110",
    "1110110010110100",
    "1110110011010111",
    "1110110111011011",
    "1110111100001001",
    "1110111111001111",
    "1111000000101011",
    "1111000011101111",
    "1111001110000100",
    "1111100100100101",
    "1111110111010101",
    "1111001010001001",
    "1110011100101010",
    "1101111000001110",
    "1101100011110100",
    "1101100001100001",
    "1101101101111111",
    "1110000010110011",
    "1110011001000110",
    "1110101100011011",
    "1110111011110010",
    "1111001000010101",
    "1111010011010010",
    "1111011100111111",
    "1111100101110100",
    "1111110000000001",
    "1111111101110001",
    "1111110000011100",
    "1111011100001001",
    "1111001000100000",
    "1110111001001011",
    "1110110001101001",
    "1110110100001011",
    "1110111111001101",
    "1111001110010001",
    "1111011100011011",
    "1111100101100111",
    "1111101000100001",
    "1111100110000100",
    "1111100000001010",
    "1111011001010110",
    "1111010011010000",
    "1111001110001010",
    "1111001001101010",
    "1111000101000001",
    "1111000000000111",
    "1110111011110010",
    "1110111011101000",
    "1111000100111011",
    "1111011010010011",
    "1111111010110101",
    "1111011110010100",
    "1110111000111010",
    "1110011100011011",
    "1110001110010010",
    "1110001111100110",
    "1110011100000100",
    "1110101100110010",
    "1110111011001010",
    "1111000101000001",
    "1111001101111000",
    "1111011010011000",
    "1111101101011010",
    "1111111001001000",
    "1111011101110111",
    "1111000111000011",
    "1110111001111111",
    "1110111000100111",
    "1110111111101100",
    "1111001001010001",
    "1111001111101100",
    "1111001111111011",
    "1111001010111000",
    "1111000011111001",
    "1110111110001101",
    "1110111101011100",
    "1111000101010011",
    "1111010111001110",
    "1111110001110001",
    "1111101111000011",
    "1111010001010111",
    "1110111010011101",
    "1110101101110000",
    "1110101100100110",
    "1110110100011111",
    "1111000000001010",
    "1111001010011000",
    "1111001110110011",
    "1111001100001100",
    "1111000100000011",
    "1110111000111100",
    "1110110000001111",
    "1110110000011111",
    "1110111100110000",
    "1111010100001011",
    "1111110001111010",
    "1111110001100011",
    "1111011100001110",
    "1111010001011110",
    "1111010001010101",
    "1111010111101101",
    "1111100000101011",
    "1111101011011111",
    "1111111001000000",
    "1111110101010111",
    "1111011111111101",
    "1111001010011011",
    "1110111001100011",
    "1110110010010000",
    "1110110111010001",
    "1111000101111011",
    "1111010111111001",
    "1111100110111111",
    "1111110000110110",
    "1111111000001000",
    "1111111110101101",
    "1111110000011110",
    "1111011101000100",
    "1111001000101000",
    "1110111001101010",
    "1110110101100010",
    "1110111101100100",
    "1111001110001010",
    "1111100001001000",
    "1111110000100111",
    "1111111001001100",
    "1111111011101110",
    "1111111101101111",
    "1111111001111100",
    "1111100111011001",
    "1111001011101111",
    "1110101101001111",
    "1110010100011000",
    "1110001000100010",
    "1110001101110011",
    "1110100010001111",
    "1110111110101000",
    "1111011011001001",
    "1111110001100110",
    "1111111111000001",
    "1111111100011101",
    "1111111111011101",
    "1111111000011111",
    "1111101111011111",
    "1111101010011010",
    "1111101101011010",
    "1111111010010010",
    "1111110000011110",
    "1111010111100010",
    "1111000000101001",
    "1110110001011001",
    "1110101101100100",
    "1110110110001000",
    "1111001001001011",
    "1111100010011001",
    "1111111100000100",
    "1111101110101110",
    "1111100001100111",
    "1111011110101001",
    "1111100110100110",
    "1111111000101111",
    "1111101101101101",
    "1111010001011111",
    "1110111000000001",
    "1110100110001110",
    "1110100001010100",
    "1110101101101110",
    "1111001011001100",
    "1111110100000011",
    "1111100000100110",
    "1110111100010110",
    "1110100110001000",
    "1110100001000101",
    "1110101011100001",
    "1110111110110011",
    "1111010010110001",
    "1111100000111101",
    "1111100101110111",
    "1111100010001010",
    "1111011000111111",
    "1111001101111011",
    "1111000101001000",
    "1111000011101001",
    "1111001101000010",
    "1111100010000011",
    "1111111111111000",
    "1111011111011110",
    "1111000010010111",
    "1110101110000101",
    "1110100110010101",
    "1110101010100011",
    "1110110110011111",
    "1111000100101111",
    "1111010000100100",
    "1111010111101100",
    "1111011010011001",
    "1111011100000101",
    "1111100010001101",
    "1111110000011000",
    "1111111001101101",
    "1111100000000111",
    "1111001001000110",
    "1110111010000111",
    "1110110110000011",
    "1110111011100001",
    "1111000101011101",
    "1111001110101000",
    "1111010011011111",
    "1111010011000000",
    "1111001110111000",
    "1111001010000100",
    "1111000111011010",
    "1111001001011000",
    "1111010001111011",
    "1111100001111000",
    "1111111000010001",
    "1111101110011010",
    "1111010111100000",
    "1111000111111100",
    "1111000010101110",
    "1111000111100000",
    "1111010001100111",
    "1111011001100111",
    "1111011000110000",
    "1111001100000010",
    "1110110101110001",
    "1110011100100011",
    "1110001000001001",
    "1101111110011100",
    "1110000001010010",
    "1110001101111111",
    "1110011111011001",
    "1110110000010111",
    "1110111101010100",
    "1111000101000000",
    "1111001000011010",
    "1111001011101111",
    "1111010100001101",
    "1111100100100010",
    "1111111100001010",
    "1111101000111010",
    "1111010000101001",
    "1110111111110001",
    "1110111001010001",
    "1110111101000000",
    "1111000111001001",
    "1111010011011100",
    "1111100000001111",
    "1111101110001110",
    "1111111110110111",
    "1111101101110111",
    "1111011001101011",
    "1111000110110111",
    "1110111000011000",
    "1110110001000011",
    "1110110001011111",
    "1110110111100111",
    "1111000001001100",
    "1111001100101000",
    "1111011001111101",
    "1111101010011111",
    "1111111110110110",
    "1111101001100001",
    "1111010000111011",
    "1110111011011101",
    "1110101100111010",
    "1110100111011011",
    "1110101011000010",
    "1110110101001011",
    "1111000001111011",
    "1111001101101001",
    "1111010110100000",
    "1111011101110101",
    "1111100110100110",
    "1111110010100011",
    "1111111110011101",
    "1111101111010000",
    "1111100100011100",
    "1111100010010101",
    "1111101011010000",
    "1111111101110101",
    "1111101010100000",
    "1111010010111110",
    "1110111111000111",
    "1110110000101100",
    "1110100111111110",
    "1110100100101001",
    "1110100110100101",
    "1110101101011001",
    "1110111000111111",
    "1111001011001110",
    "1111100101110001",
    "1111110111111011",
    "1111010000110101",
    "1110101010011101",
    "1110001010111101",
    "1101110110110100",
    "1101110000101011",
    "1101110111100011",
    "1110000110111110",
    "1110011011100011",
    "1110110100110111",
    "1111010011011010",
    "1111110111010101",
    "1111100010000000",
    "1110111101111111",
    "1110100001100111",
    "1110010001000010",
    "1110001101111011",
    "1110010101011010",
    "1110100010010010",
    "1110101111000101",
    "1110110111111010",
    "1110111110110110",
    "1111001010001111",
    "1111011111000100",
    "1111111110010101",
    "1111011100110101",
    "1110111011110101",
    "1110100110100100",
    "1110100010000010",
    "1110101101100110",
    "1111000010010000",
    "1111010110111100",
    "1111100101010000",
    "1111101101101001",
    "1111110110011000",
    "1111111011010001",
    "1111100110001000",
    "1111001101001110",
    "1110110111010000",
    "1110101011000111",
    "1110101101001110",
    "1110111100110111",
    "1111010011100100",
    "1111101011001001",
    "1111111110101101",
    "1111101001011111",
    "1111010010111001",
    "1110111011000100",
    "1110100101101001",
    "1110010111000100",
    "1110010100000001",
    "1110011110000101",
    "1110110001100110",
    "1111001000000100",
    "1111011010111101",
    "1111101000001011",
    "1111110011111001",
    "1111111100000000",
    "1111100011111011",
    "1111000101000101",
    "1110100110101000",
    "1110010001101110",
    "1110001101010110",
    "1110011011100101",
    "1110110111010110",
    "1111010111011111",
    "1111110010100100",
    "1111111101011101",
    "1111111000110010",
    "1111111011010011",
    "1111111111101101",
    "1111111100000101",
    "1111111011000001",
    "1111111011011001",
    "1111111011011010",
    "1111111001001011",
    "1111110100110001",
    "1111110010011111",
    "1111110111111100",
    "1111110111111111",
    "1111011110110101",
    "1111000010100001",
    "1110101010011000",
    "1110011011111111",
    "1110011010000010",
    "1110100010111110",
    "1110110001011111",
    "1111000000000000",
    "1111001001111111",
    "1111001110000111",
    "1111010000101110",
    "1111011000011101",
    "1111101001111010",
    "1111111010001110",
    "1111011000110111",
    "1110111001110000",
    "1110100011111000",
    "1110011100000100",
    "1110100001111110",
    "1110101111110110",
    "1110111111000000",
    "1111001010011011",
    "1111010000001111",
    "1111010001111101",
    "1111010001010100",
    "1111010001000000",
    "1111010110010000",
    "1111100100110011",
    "1111111100110111",
    "1111100100100100",
    "1111000110000100",
    "1110101110000100",
    "1110100000101100",
    "1110100000000111",
    "1110101010010011",
    "1110111001111010",
    "1111001001010101",
    "1111010011100100",
    "1111010110011101",
    "1111010011000101",
    "1111001011100110",
    "1111000011001010",
    "1110111100011001",
    "1110111000110100",
    "1110111011010110",
    "1111000110110001",
    "1111011011101000",
    "1111111000010100",
    "1111100111101100",
    "1111001010101000",
    "1110110110001000",
    "1110101110010110",
    "1110110010011111",
    "1110111101101000",
    "1111001100111000",
    "1111011111111000",
    "1111110110101110",
    "1111101110111101",
    "1111010100100100",
    "1110111110011100",
    "1110110000000111",
    "1110101100100011",
    "1110110011011100",
    "1111000011000101",
    "1111011010011000",
    "1111110110110011",
    "1111101011000001",
    "1111001110111101",
    "1110111001001110",
    "1110101100101101",
    "1110101010110101",
    "1110110011011000",
    "1111000010110001",
    "1111010100100100",
    "1111100110111110",
    "1111111010011011",
    "1111110000001111",
    "1111011001000010",
    "1111000001010100",
    "1110101010111010",
    "1110011001000001",
    "1110001111110011",
    "1110010001100001",
    "1110011110111010",
    "1110111000000110",
    "1111011011100011",
    "1111111001011011",
    "1111001010100010",
    "1110011101100001",
    "1101111000110000",
    "1101100001011001",
    "1101011010000111",
    "1101100001001111",
    "1101110010000110",
    "1110000111011000",
    "1110011100000001",
    "1110101101010010",
    "1110111010110111",
    "1111000101100101",
    "1111001111100110",
    "1111011010010011",
    "1111100100011101",
    "1111101011110011",
    "1111101101111100",
    "1111101001101001",
    "1111100000001000",
    "1111010011110100",
    "1111000111111001",
    "1110111111011100",
    "1110111011110111",
    "1110111110111010",
    "1111001010011110",
    "1111011110110101",
    "1111111010100101",
    "1111100110000000",
    "1111001000011110",
    "1110110001010111",
    "1110100011111011",
    "1110100000101011",
    "1110100100011010",
    "1110101010100101",
    "1110101111010001",
    "1110110000001100",
    "1110110000000101",
    "1110110101010000",
    "1111000101001000",
    "1111100001111011",
    "1111111000010100",
    "1111010010110011",
    "1110110110101100",
    "1110101010110100",
    "1110110000011111",
    "1111000010010101",
    "1111011000001000",
    "1111101010100100",
    "1111110111100010",
    "1111111100111000",
    "1111101110000010",
    "1111011001111010",
    "1111000001110011",
    "1110101011100000",
    "1110011110010100",
    "1110100000000000",
    "1110110011001010",
    "1111010100000110",
    "1111111010101111",
    "1111100001100110",
    "1111000111010110",
    "1110111000010110",
    "1110110011000011",
    "1110110101001000",
    "1110111011101111",
    "1111000101001000",
    "1111010001100110",
    "1111100001101011",
    "1111110100010110",
    "1111111001011001",
    "1111101100010111",
    "1111101000010010",
    "1111101101111001",
    "1111111010101111",
    "1111110101100001",
    "1111100111101000",
    "1111011110001010",
    "1111011001111010",
    "1111011011101101",
    "1111100100011000",
    "1111110011111110",
    "1111110110011110",
    "1111011110001111",
    "1111001000000100",
    "1110111000101100",
    "1110110011101100",
    "1110111000111100",
    "1111000011101110",
    "1111001110111101",
    "1111011001000111",
    "1111100011100010",
    "1111110000101000",
    "1111111110011000",
    "1111101010111101",
    "1111011000000011",
    "1111001010001111",
    "1111000110000011",
    "1111001100001110",
    "1111011001011001",
    "1111100111111101",
    "1111110011010111",
    "1111111100101001",
    "1111110111101000",
    "1111100101101100",
    "1111001100011110",
    "1110101111100001",
    "1110010101100101",
    "1110000101101100",
    "1110000100111011",
    "1110010011001111",
    "1110101011100001",
    "1111000110011010",
    "1111011101100001",
    "1111110000011111",
    "1111111100111101",
    "1111101000000111",
    "1111010000011110",
    "1110111000111110",
    "1110100111000001",
    "1110011111110101",
    "1110100110100101",
    "1110111001110111",
    "1111010011011010",
    "1111101011110000",
    "1111111100111100",
    "1111111010111000",
    "1111111001111010",
    "1111111101101000",
    "1111111100011000",
    "1111110110000100",
    "1111101111101101",
    "1111101001111101",
    "1111100111100001",
    "1111101011010101",
    "1111110110110101",
    "1111110110111101",
    "1111100001111101",
    "1111001111100011",
    "1111000100110001",
    "1111000100001000",
    "1111001011110111",
    "1111010111000100",
    "1111100001100100",
    "1111101001011011",
    "1111101111010110",
    "1111110101100101",
    "1111111110010000",
    "1111110101101011",
    "1111100111100011",
    "1111011010101000",
    "1111010001111110",
    "1111001110011111",
    "1111001110111011",
    "1111010000111001",
    "1111010001111001",
    "1111010000111001",
    "1111001110100001",
    "1111001101100000",
    "1111010011001111",
    "1111100100010111",
    "1111111110101000",
    "1111011001100111",
    "1110110100101001",
    "1110011010101011",
    "1110010101010011",
    "1110101001000110",
    "1111010010101110",
    "1111111000101101",
    "1111000110110100",
    "1110100011001010",
    "1110010100001000",
    "1110011000010110",
    "1110101010011000",
    "1111000101100101",
    "1111100110011101",
    "1111110101001011",
    "1111001111010110",
    "1110101100000111",
    "1110001111110101",
    "1101111110100001",
    "1101111011011000",
    "1110000101001101",
    "1110010110011010",
    "1110101000011011",
    "1110110101101010",
    "1110111101001001",
    "1111000100001000",
    "1111010001001010",
    "1111101001000010",
    "1111110100000110",
    "1111001100110010",
    "1110101001101101",
    "1110010010100110",
    "1110001100001001",
    "1110010100100100",
    "1110100101100000",
    "1110111000010001",
    "1111001000100000",
    "1111010111100111",
    "1111101010001000",
    "1111111101010111",
    "1111011111100001",
    "1111000001001000",
    "1110101010000110",
    "1110100000111101",
    "1110101001011001",
    "1111000010001000",
    "1111100100001010",
    "1111111000111011",
    "1111011011111010",
    "1111000111110111",
    "1110111100011001",
    "1110111000010110",
    "1110111010101111",
    "1111000011000110",
    "1111010010111110",
    "1111101011001111",
    "1111110110001100",
    "1111010101110100",
    "1110111001011101",
    "1110100110111111",
    "1110100010001111",
    "1110101100000111",
    "1111000010000110",
    "1111011111011010",
    "1111111111100101",
    "1111100001011110",
    "1111000111010011",
    "1110110100000110",
    "1110101001000111",
    "1110100101111011",
    "1110101000101111",
    "1110101111100011",
    "1110110111110010",
    "1111000001100111",
    "1111010000100011",
    "1111100111100000",
    "1111111000111110",
    "1111010100001101",
    "1110110000110011",
    "1110010101011111",
    "1110000111110010",
    "1110001010000001",
    "1110011000110010",
    "1110101110010001",
    "1111000111000110",
    "1111100010100001",
    "1111111110111100",
    "1111011101110011",
    "1110111101011011",
    "1110100010101100",
    "1110010010111000",
    "1110010010010000",
    "1110100000100011",
    "1110111000100111",
    "1111010011100100",
    "1111101010011100",
    "1111111001111001",
    "1111111011011001",
    "1111110000110100",
    "1111100010111011",
    "1111010001011010",
    "1111000000001100",
    "1110110100000011",
    "1110110000011111",
    "1110110110110110",
    "1111000100011100",
    "1111010100010010",
    "1111100001111000",
    "1111101010110110",
    "1111101111101111",
    "1111110010100100",
    "1111110100001100",
    "1111110100100010",
    "1111110011101000",
    "1111110011010001",
    "1111110110101010",
    "1111111111101011",
    "1111110010011000",
    "1111100011000001",
    "1111010111110111",
    "1111010110100000",
    "1111100010001011",
    "1111111000110110",
    "1111101101101000",
    "1111011011011101",
    "1111011000010000",
    "1111100110001101",
    "1111111111000101",
    "1111100000010010",
    "1111000110100111",
    "1110111000100111",
    "1110110111101111",
    "1111000000101100",
    "1111001101100001",
    "1111011000100111",
    "1111011110110110",
    "1111100000010010",
    "1111011110101110",
    "1111011011111101",
    "1111011000100011",
    "1111010101010101",
    "1111010101001011",
    "1111011011001010",
    "1111101000111110",
    "1111111110001011",
    "1111101000100101",
    "1111010000101011",
    "1110111111011110",
    "1110111000101100",
    "1110111100000101",
    "1111000111111110",
    "1111011011100101",
    "1111110101010011",
    "1111101101010001",
    "1111001111110011",
    "1110110111001101",
    "1110100111001101",
    "1110100010000101",
    "1110101000001001",
    "1110110101100111",
    "1111000101010011",
    "1111010010010010",
    "1111011001110101",
    "1111011111010010",
    "1111101000100101",
    "1111111010001001",
    "1111101010101000",
    "1111001010010001",
    "1110101100100110",
    "1110011000111100",
    "1110010011111001",
    "1110011100011011",
    "1110101100010011",
    "1110111100010110",
    "1111000111010001",
    "1111001011101101",
    "1111001100000101",
    "1111001011001111",
    "1111001100010001",
    "1111010100000001",
    "1111100101100111",
    "1111111111100011",
    "1111011111011010",
    "1111000001001010",
    "1110101011100011",
    "1110100010011101",
    "1110100111000001",
    "1110110110010010",
    "1111001001110101",
    "1111011011010011",
    "1111100101100100",
    "1111100110100101",
    "1111100000100111",
    "1111011000100010",
    "1111010100001011",
    "1111010111101111",
    "1111100010011100",
    "1111101111000110",
    "1111110110110010",
    "1111110011101111",
    "1111100100110110",
    "1111001110011100",
    "1110111000101000",
    "1110101101011001",
    "1110110100001000",
    "1111001110011011",
    "1111110111110011",
    "1111011000111111",
    "1110101110111011",
    "1110010010000000",
    "1110000101011010",
    "1110000110101111",
    "1110001111101000",
    "1110011001110111",
    "1110100001000101",
    "1110100101000110",
    "1110101011001100",
    "1110111001010000",
    "1111010001111000",
    "1111110011011100",
    "1111101000100110",
    "1111001010000111",
    "1110110111001001",
    "1110110010111000",
    "1110111010101010",
    "1111000111110111",
    "1111010011100100",
    "1111011001011110",
    "1111011100001001",
    "1111100010001101",
    "1111110000101010",
    "1111110110110011",
    "1111010111111001",
    "1110111010100000",
    "1110100110011011",
    "1110100001000101",
    "1110101010100010",
    "1110111101000100",
    "1111010000111001",
    "1111011111001100",
    "1111100100101001",
    "1111100010011010",
    "1111011011100001",
    "1111010011011000",
    "1111001110001010",
    "1111001111110110",
    "1111011010101000",
    "1111101101111110",
    "1111111001010100",
    "1111100000001100",
    "1111001011010001",
    "1110111110011011",
    "1110111011110000",
    "1111000010000000",
    "1111001101000100",
    "1111011000010011",
    "1111011111110000",
    "1111100001101110",
    "1111011110100110",
    "1111010111011010",
    "1111001110001100",
    "1111000100101010",
    "1110111011011000",
    "1110110010010000",
    "1110101001010000",
    "1110100001001101",
    "1110011100100101",
    "1110011101010110",
    "1110100011110110",
    "1110101110010110",
    "1110111001111101",
    "1111000100001101",
    "1111001011100000",
    "1111001111011010",
    "1111010001010100",
    "1111010011010111",
    "1111011000011110",
    "1111100100100100",
    "1111111001110110",
    "1111101000100100",
    "1111000110001101",
    "1110100100110100",
    "1110001010010100",
    "1101111010111100",
    "1101111000100101",
    "1110000000110000",
    "1110001111110000",
    "1110100100101110",
    "1110111111100100",
    "1111011111111101",
    "1111111011101110",
    "1111011000000001",
    "1110111001111010",
    "1110100110000110",
    "1110100000011111",
    "1110101001110111",
    "1111000000010100",
    "1111011111101011",
    "1111111110111001",
    "1111100010101110",
    "1111010010000110",
    "1111010001011001",
    "1111100000011100",
    "1111111010111011",
    "1111100110110101",
    "1111001101111000",
    "1111000000010101",
    "1110111111101110",
    "1111001001001011",
    "1111010110101101",
    "1111100001110001",
    "1111100101100000",
    "1111100010010111",
    "1111011111000101",
    "1111100011101010",
    "1111110100101110",
    "1111101110010111",
    "1111001011110000",
    "1110101011100001",
    "1110010100100101",
    "1110001010001110",
    "1110001010100110",
    "1110010000111011",
    "1110011000100101",
    "1110011110110001",
    "1110100011110110",
    "1110101011111101",
    "1110111100110111",
    "1111011001110100",
    "1111111110010011",
    "1111010001111011",
    "1110101010001111",
    "1110001111001111",
    "1110000101110100",
    "1110001101101001",
    "1110100000110110",
    "1110110111111001",
    "1111001100101110",
    "1111011011111101",
    "1111100101000011",
    "1111101001101111",
    "1111101110111011",
    "1111111010100001",
    "1111110000101000",
    "1111010011111011",
    "1110110100011111",
    "1110011001001100",
    "1110000111111111",
    "1110000011101100",
    "1110001100010001",
    "1110100000100110",
    "1110111110010100",
    "1111100001001101",
    "1111111100000100",
    "1111011111100011",
    "1111001101111111",
    "1111001001101010",
    "1111010001111110",
    "1111100011000011",
    "1111110111100101",
    "1111110010101010",
    "1111011011001110",
    "1111000001001000",
    "1110100101001101",
    "1110001011100011",
    "1101111001010011",
    "1101110010100010",
    "1101111010011001",
    "1110010000000111",
    "1110101110000101",
    "1111001100110011",
    "1111100101000001",
    "1111110010110110",
    "1111110110110101",
    "1111110101011001",
    "1111110110001111",
    "1111111111111001",
    "1111101011011111",
    "1111001111110110",
    "1110110100000011",
    "1110011111111011",
    "1110011000110100",
    "1110100000001111",
    "1110110011000110",
    "1111001011010011",
    "1111100010111001",
    "1111110101100100",
    "1111111110010101",
    "1111111000011011",
    "1111110111100010",
    "1111111010010101",
    "1111111111000101",
    "1111111100100111",
    "1111111011101001",
    "1111111111101110",
    "1111110101000111",
    "1111100110011110",
    "1111010111101010",
    "1111001101001010",
    "1111001010100101",
    "1111010000101100",
    "1111011101001001",
    "1111101011010110",
    "1111110110111100",
    "1111111100111101",
    "1111111101011101",
    "1111111100101011",
    "1111111111100010",
    "1111110011111100",
    "1111100001010101",
    "1111001100100011",
    "1110111011110010",
    "1110110100001000",
    "1110110111111111",
    "1111000101001101",
    "1111010110000001",
    "1111100100100111",
    "1111101110010001",
    "1111110101010111",
    "1111111110101000",
    "1111110010110011",
    "1111011110100001",
    "1111000111010000",
    "1110110010001000",
    "1110100100001010",
    "1110100000000010",
    "1110100100100101",
    "1110101101110011",
    "1110110111100111",
    "1110111111011111",
    "1111000110011010",
    "1111010000110101",
    "1111100010100001",
    "1111111100000010",
    "1111100101011111",
    "1111000111111111",
    "1110110001100111",
    "1110100110011010",
    "1110100111100111",
    "1110110010001101",
    "1111000000010100",
    "1111001100101110",
    "1111010100000110",
    "1111010110100100",
    "1111011000101100",
    "1111011111101011",
    "1111101110101010",
    "1111111010101001",
    "1111100001100110",
    "1111001101000000",
    "1111000011100110",
    "1111001100000100",
    "1111101000001011",
    "1111101100111001",
    "1110111011110111",
    "1110001111100011",
    "1101110001000111",
    "1101100101010010",
    "1101101100100000",
    "1110000010011101",
    "1110100001110000",
    "1111000110011101",
    "1111101100101110",
    "1111101110011100",
    "1111001110010001",
    "1110110110000001",
    "1110100111111001",
    "1110100100110001",
    "1110101011000100",
    "1110110110011010",
    "1111000010100001",
    "1111001100001001",
    "1111010010011010",
    "1111011000010101",
    "1111100000100111",
    "1111101011010110",
    "1111110110001001",
    "1111111100111101",
    "1111111100101110",
    "1111110100111011",
    "1111101000101010",
    "1111100000010001",
    "1111100100101001",
    "1111111001000000",
    "1111100110110111",
    "1111000100110111",
    "1110101011100011",
    "1110100001011110",
    "1110100111101100",
    "1110111001000110",
    "1111001100111100",
    "1111011011110000",
    "1111100001111110",
    "1111100000010001",
    "1111011010101000",
    "1111010101110010",
    "1111010110101000",
    "1111100000111001",
    "1111110100110001",
    "1111101111111001",
    "1111010001000111",
    "1110110100010000",
    "1110011110001010",
    "1110010010010100",
    "1110010010011010",
    "1110011100111111",
    "1110101110100011",
    "1111000010110011",
    "1111010101011000",
    "1111100011011101",
    "1111101100000011",
    "1111101110111100",
    "1111101110010001",
    "1111101111001100",
    "1111110111000111",
    "1111110110110011",
    "1111011011100011",
    "1110111100111111",
    "1110100010101001",
    "1110010010100100",
    "1110010000001111",
    "1110011010100000",
    "1110101011110101",
    "1110111101110111",
    "1111001011001110",
    "1111010001111110",
    "1111010011101110",
    "1111010010011001",
    "1111010000101001",
    "1111010010101100",
    "1111011010111010",
    "1111101001011001",
    "1111111100001011",
    "1111110000110000",
    "1111100001001010",
    "1111010111100000",
    "1111010100111011",
    "1111010111100111",
    "1111011100010001",
    "1111011111100100",
    "1111011110101101",
    "1111011000101100",
    "1111001110110110",
    "1111000011011111",
    "1110111001011101",
    "1110110011001010",
    "1110110001010010",
    "1110110011111001",
    "1110111010001011",
    "1111000010010000",
    "1111001010011110",
    "1111010001100111",
    "1111010111001001",
    "1111011010110010",
    "1111011101011100",
    "1111100010101110",
    "1111101111011100",
    "1111111010010010",
    "1111011100010111",
    "1110111011111111",
    "1110011111111011",
    "1110001101101001",
    "1110001000010011",
    "1110010000011001",
    "1110100011101110",
    "1110111110101001",
    "1111011100111000",
    "1111111010010111",
    "1111101100010001",
    "1111011010000110",
    "1111010001001111",
    "1111010010001000",
    "1111011011110111",
    "1111101100100011",
    "1111111110110000",
    "1111101001101101",
    "1111010111101101",
    "1111001011100000",
    "1111000110000000",
    "1111000101110110",
    "1111001000000100",
    "1111001001100011",
    "1111001000011010",
    "1111000100011010",
    "1110111110100110",
    "1110111000011101",
    "1110110100010111",
    "1110110110100010",
    "1111000010101011",
    "1111011001001011",
    "1111110110100110",
    "1111101011100011",
    "1111010100010111",
    "1111001000111111",
    "1111001011111100",
    "1111011010110111",
    "1111101111011000",
    "1111111011011100",
    "1111100110111000",
    "1111010010010101",
    "1110111101000010",
    "1110101000010011",
    "1110010111100010",
    "1110001110010111",
    "1110010000101001",
    "1110011111111010",
    "1110111000101100",
    "1111010100110011",
    "1111101101001011",
    "1111111100111001",
    "1111111001110010",
    "1111110000010110",
    "1111100001010100",
    "1111001010100110",
    "1110110000000011",
    "1110011001001011",
    "1110001100100101",
    "1110001110100011",
    "1110011101111111",
    "1110110100001011",
    "1111001001101010",
    "1111011000110000",
    "1111100000000111",
    "1111100010001000",
    "1111100010000101",
    "1111100101000001",
    "1111110000000000",
    "1111111100001101",
    "1111100010111000",
    "1111001001111100",
    "1110111000000011",
    "1110110000111001",
    "1110110101000000",
    "1111000001000111",
    "1111001111011110",
    "1111011010111111",
    "1111100000000101",
    "1111011101101001",
    "1111010101110111",
    "1111001100011001",
    "1111000101000011",
    "1111000011100110",
    "1111001010000111",
    "1111011000110010",
    "1111101101110110",
    "1111111010100011",
    "1111100101011011",
    "1111010110111100",
    "1111010001011001",
    "1111010100101111",
    "1111011110010100",
    "1111101001011110",
    "1111110000001101",
    "1111101101101100",
    "1111100000111101",
    "1111001101000100",
    "1110110111011000",
    "1110100101010101",
    "1110011010001111",
    "1110011000110000",
    "1110100010111001",
    "1110110111111001",
    "1111010100011111",
    "1111110011111011",
    "1111101111001010",
    "1111011000110111",
    "1111001011110101",
    "1111001000110111",
    "1111001101101000",
    "1111010110001000",
    "1111011110110001",
    "1111100100101111",
    "1111100111001000",
    "1111100110010000",
    "1111100011000011",
    "1111011111011010",
    "1111011101001111",
    "1111011110000010",
    "1111100011110011",
    "1111101111100011",
    "1111111110110111",
    "1111101000100000",
    "1111001111111111",
    "1110111001011101",
    "1110101001000110",
    "1110100001101011",
    "1110100010111110",
    "1110101010010001",
    "1110110100001101",
    "1110111101100000",
    "1111000011110110",
    "1111000110111100",
    "1111001000100000",
    "1111001011101101",
    "1111010010011101",
    "1111011011101101",
    "1111100100010000",
    "1111101000011111",
    "1111100110000110",
    "1111011101111111",
    "1111010100110111",
    "1111010001100010",
    "1111011001000111",
    "1111101100010001",
    "1111111000110010",
    "1111011100101101",
    "1111000101110111",
    "1110111000011000",
    "1110110101000000",
    "1110111001011000",
    "1111000001101001",
    "1111001010010100",
    "1111010000111101",
    "1111010100100000",
    "1111010101011000",
    "1111010100110111",
    "1111010100101110",
    "1111010110011000",
    "1111011010100110",
    "1111100001111101",
    "1111101101000110",
    "1111111100100100",
    "1111110000001110",
    "1111011011010110",
    "1111000111100111",
    "1110110111011111",
    "1110101100011011",
    "1110100110110001",
    "1110100101101100",
    "1110101000011011",
    "1110110000000111",
    "1110111111000100",
    "1111010110011000",
    "1111110100101100",
    "1111101010110100",
    "1111001110111011",
    "1110111101001010",
    "1110111000101010",
    "1110111111111010",
    "1111001101000111",
    "1111011001100101",
    "1111100000001100",
    "1111100001101011",
    "1111100100110001",
    "1111110000100010",
    "1111110111000010",
    "1111010011110100",
    "1110101101101101",
    "1110001110010100",
    "1101111101100000",
    "1101111110000100",
    "1110001101010110",
    "1110100111100101",
    "1111001000011110",
    "1111101011110111",
    "1111110001000110",
    "1111010010000110",
    "1110111010110010",
    "1110101101101001",
    "1110101100001110",
    "1110110100111110",
    "1111000011100100",
    "1111010101000001",
    "1111101001100101",
    "1111111101100100",
    "1111100000011100",
    "1111000001011111",
    "1110100101000011",
    "1110010000001010",
    "1110000111110010",
    "1110001110100100",
    "1110100001110000",
    "1110111011000001",
    "1111010011001000",
    "1111100100001011",
    "1111101110111001",
    "1111111001011111",
    "1111110110010101",
    "1111011101100110",
    "1110111110101011",
    "1110100000111011",
    "1110001011110111",
    "1110000101100111",
    "1110001111101011",
    "1110100101010000",
    "1110111110110110",
    "1111010110110001",
    "1111101100100100",
    "1111111011110111",
    "1111011111011111",
    "1110111110010100",
    "1110011011111101",
    "1101111111010111",
    "1101101111110001",
    "1101110010011111",
    "1110001001010001",
    "1110110000100100",
    "1111100000111011",
    "1111101110011000",
    "1111000101010111",
    "1110101000110100",
    "1110011011000111",
    "1110011100001110",
    "1110101000101101",
    "1110111011010011",
    "1111001110101101",
    "1111011110101101",
    "1111101000110100",
    "1111101101011000",
    "1111110000001100",
    "1111110111000111",
    "1111111001010010",
    "1111100000101100",
    "1111000011110100",
    "1110101010011110",
    "1110011100000001",
    "1110011100011110",
    "1110101010100000",
    "1111000000000011",
    "1111010110010000",
    "1111100111001001",
    "1111110001000000",
    "1111111000011000",
    "1111111100011001",
    "1111101001011100",
    "1111001111001000",
    "1110110011010010",
    "1110011101110111",
    "1110010101011011",
    "1110011101001010",
    "1110110010000010",
    "1111001101011011",
    "1111101001010010",
    "1111111110110001",
    "1111101100001101",
    "1111011110011111",
    "1111010101111100",
    "1111010011001111",
    "1111010111000011",
    "1111100001100001",
    "1111110000000010",
    "1111111110101110",
    "1111110110001011",
    "1111110010000111",
    "1111110110010011",
    "1111111110101110",
    "1111110001000010",
    "1111100101100010",
    "1111011111011010",
    "1111011111001010",
    "1111100011001000",
    "1111101000001100",
    "1111101100000011",
    "1111101110100000",
    "1111110000100111",
    "1111110011110010",
    "1111111001001100",
    "1111111111001001",
    "1111110110000011",
    "1111101100010010",
    "1111100010111011",
    "1111011011000100",
    "1111010110000001",
    "1111010101000110",
    "1111011000010110",
    "1111011110000101",
    "1111100011001111",
    "1111100100100100",
    "1111100000010111",
    "1111010110111110",
    "1111001010110000",
    "1110111111111010",
    "1110111010000100",
    "1110111011011001",
    "1111000110000100",
    "1111011010100101",
    "1111110110110011",
    "1111101001010011",
    "1111001011011000",
    "1110110100011101",
    "1110100111100101",
    "1110100101110001",
    "1110101100101101",
    "1110110111001001",
    "1111000000101110",
    "1111001001010110",
    "1111010100100010",
    "1111100110001101",
    "1111111111100001",
    "1111100010010100",
    "1111000100110100",
    "1110101110101001",
    "1110100101001101",
    "1110101001000111",
    "1110110110001011",
    "1111000101101111",
    "1111010001011100",
    "1111010101101111",
    "1111010011010111",
    "1111001100111111",
    "1111000101110110",
    "1111000000010100",
    "1110111100011011",
    "1110111000111010",
    "1110110100010101",
    "1110101101110000",
    "1110100101100101",
    "1110011101101001",
    "1110010111111100",
    "1110010110111111",
    "1110011110011011",
    "1110110000011110",
    "1111001101000100",
    "1111110001000111",
    "1111101001100111",
    "1111001001110100",
    "1110110100011111",
    "1110101011111100",
    "1110101101110101",
    "1110110101000011",
    "1110111100100011",
    "1111000000010101",
    "1110111111011111",
    "1110111011101010",
    "1110110110110111",
    "1110110100101111",
    "1110111010100010",
    "1111001011100000",
    "1111100111101000",
    "1111110100111100",
    "1111010001100001",
    "1110110101000011",
    "1110100100010000",
    "1110100000111001",
    "1110101000101010",
    "1110110111100000",
    "1111001011001100",
    "1111100010010000",
    "1111111011111011",
    "1111101001010101",
    "1111010001001100",
    "1110111111000101",
    "1110110101110110",
    "1110110111001000",
    "1111000000111011",
    "1111001110010110",
    "1111011010000001",
    "1111011111011111",
    "1111011101000111",
    "1111010100010111",
    "1111001000101100",
    "1110111110000100",
    "1110110111001001",
    "1110110100010000",
    "1110110100000001",
    "1110110100110011",
    "1110110110110010",
    "1110111100110011",
    "1111001001010101",
    "1111011100011011",
    "1111110011000101",
    "1111110111111000",
    "1111101001010000",
    "1111100011110001",
    "1111100111000011",
    "1111101110111010",
    "1111110101101010",
    "1111110110110001",
    "1111110000011110",
    "1111100100011101",
    "1111010110101100",
    "1111001011100011",
    "1111000110011011",
    "1111001000100101",
    "1111010000100111",
    "1111011011111101",
    "1111101000000100",
    "1111110010110100",
    "1111111010101011",
    "1111111110000100",
    "1111111011001111",
    "1111110001001010",
    "1111100000110011",
    "1111001101000000",
    "1110111001110101",
    "1110101011001100",
    "1110100100000000",
    "1110100101010011",
    "1110101110001111",
    "1110111101010110",
    "1111010001011110",
    "1111101001110100",
    "1111111010101100",
    "1111011110010110",
    "1111000100000101",
    "1110101111000000",
    "1110100001110100",
    "1110011110011110",
    "1110100110101000",
    "1110111011001111",
    "1111011010101011",
    "1111111110111011",
    "1111010111011101",
    "1110110101010011",
    "1110011101011011",
    "1110010010011010",
    "1110010011100100",
    "1110011100100001",
    "1110101000010000",
    "1110110101010000",
    "1111000101011101",
    "1111011011101101",
    "1111111001100001",
    "1111100011010111",
    "1111000000000111",
    "1110100010111000",
    "1110010001011010",
    "1110001101101110",
    "1110010111001001",
    "1110101100110011",
    "1111001011101011",
    "1111101111100011",
    "1111101011111101",
    "1111001100001010",
    "1110110101001101",
    "1110101010000001",
    "1110101011110010",
    "1110110111110001",
    "1111001000111100",
    "1111011010111000",
    "1111101001111000",
    "1111110100101001",
    "1111111101011111",
    "1111110110110110",
    "1111100100010111",
    "1111001010110010",
    "1110101110111101",
    "1110011000011011",
    "1110001101110101",
    "1110010011000101",
    "1110100111000011",
    "1111000011010010",
    "1111011111111111",
    "1111110110100101",
    "1111111100110000",
    "1111111001111100",
    "1111111110101011",
    "1111111001100000",
    "1111110101111100",
    "1111111011101011",
    "1111110100100100",
    "1111011110010111",
    "1111001000110100",
    "1110111010100101",
    "1110110111110010",
    "1111000001100001",
    "1111010011111001",
    "1111101000011111",
    "1111111001011101",
    "1111111101110011",
    "1111111110010011",
    "1111111001110100",
    "1111101111000100",
    "1111101001011010",
    "1111101111001101",
    "1111111110101111",
    "1111100100010010",
    "1111001000011101",
    "1110110010011111",
    "1110100110111001",
    "1110100110101111",
    "1110101110100001",
    "1110111000100000",
    "1111000000011001",
    "1111000011010111",
    "1111000001100010",
    "1110111111110110",
    "1111000101011111",
    "1111010111011101",
    "1111110110010110",
    "1111100011000101",
    "1110111101011100",
    "1110100000100111",
    "1110010010011010",
    "1110010011111000",
    "1110100000011001",
    "1110110001011110",
    "1111000001111011",
    "1111001110111111",
    "1111011000110100",
    "1111011111110001",
    "1111100100001010",
    "1111100110011011",
    "1111100110000100",
    "1111100010011101",
    "1111011011100110",
    "1111010010011100",
    "1111001010111111",
    "1111001011010011",
    "1111010111011011",
    "1111101111101110",
    "1111110000000100",
    "1111001111000111",
    "1110110011111000",
    "1110100011001000",
    "1110011110011110",
    "1110100011011000",
    "1110101101010001",
    "1110110111100101",
    "1110111110101001",
    "1111000001010111",
    "1111000000111101",
    "1111000000011100",
    "1111000100011010",
    "1111010000010100",
    "1111100100100000",
    "1111111110000101",
    "1111101000010000",
    "1111010011100100",
    "1111000110101101",
    "1111000010011100",
    "1111000110000001",
    "1111010000000000",
    "1111011110101001",
    "1111101111110100",
    "1111111110010010",
    "1111101101000001",
    "1111011101010111",
    "1111010000010111",
    "1111000111001001",
    "1111000010100111",
    "1111000011001011",
    "1111001000100000",
    "1111010001010010",
    "1111011100010001",
    "1111101001011111",
    "1111111001001110",
    "1111110100101110",
    "1111100001011111",
    "1111001111110011",
    "1111000011010000",
    "1111000000000010",
    "1111001011001111",
    "1111100110101110",
    "1111110000100110",
    "1111000001010111",
    "1110010100111011",
    "1101110100001000",
    "1101100100101001",
    "1101101000001110",
    "1101111010110000",
    "1110010100001011",
    "1110101111010010",
    "1111001011011001",
    "1111101010001111",
    "1111110010101001",
    "1111001101000010",
    "1110101001100000",
    "1110001101000010",
    "1101111100100000",
    "1101111001111001",
    "1110000010010100",
    "1110010000111110",
    "1110100000110001",
    "1110101110011100",
    "1110111100011110",
    "1111001111100001",
    "1111101010011111",
    "1111110010110010",
    "1111001101111111",
    "1110101111011001",
    "1110011101100001",
    "1110011011111100",
    "1110101000100101",
    "1110111100001010",
    "1111001111000111",
    "1111011011111101",
    "1111100001010111",
    "1111100011010011",
    "1111101000001111",
    "1111110101001001",
    "1111110100001101",
    "1111010111011101",
    "1110111011110010",
    "1110101000001000",
    "1110100001010100",
    "1110100111100111",
    "1110110101110001",
    "1111000100110011",
    "1111001111010001",
    "1111010010100110",
    "1111010001010101",
    "1111010001011010",
    "1111010111101100",
    "1111100110101110",
    "1111111100110000",
    "1111101011110111",
    "1111011001000111",
    "1111010000000101",
    "1111010011010000",
    "1111100010010101",
    "1111111100001011",
    "1111100010001111",
    "1110111101101110",
    "1110011011111101",
    "1110000011010000",
    "1101111000100101",
    "1101111101100100",
    "1110010000000000",
    "1110101001111010",
    "1111000011010101",
    "1111010110111001",
    "1111100101100100",
    "1111110100011100",
    "1111111000000010",
    "1111011110100011",
    "1111000001100110",
    "1110100111000011",
    "1110010101011000",
    "1110010001011001",
    "1110011010101101",
    "1110101011111000",
    "1110111101110011",
    "1111001001110101",
    "1111001110111101",
    "1111010011101010",
    "1111100000000010",
    "1111111001010011",
    "1111100000110110",
    "1110110101111100",
    "1110010000001111",
    "1101111001000111",
    "1101110110000011",
    "1110000100110100",
    "1110011101010110",
    "1110110111010101",
    "1111001101111101",
    "1111100000111110",
    "1111110010000011",
    "1111111111001011",
    "1111110101010000",
    "1111110011001100",
    "1111111011100011",
    "1111110001111100",
    "1111011001101101",
    "1111000010101100",
    "1110110011101110",
    "1110110000011110",
    "1110110111101000",
    "1111000100011100",
    "1111010001101011",
    "1111011011110010",
    "1111100010000011",
    "1111100101100100",
    "1111101001110000",
    "1111110100000100",
    "1111110111111111",
    "1111011011000110",
    "1110111001011001",
    "1110011001110000",
    "1110000010011100",
    "1101110111101000",
    "1101111011010110",
    "1110001011011110",
    "1110100011000110",
    "1110111100100101",
    "1111010010011101",
    "1111100100000011",
    "1111110101001110",
    "1111110110100011",
    "1111011101111000",
    "1111000010101111",
    "1110101011000110",
    "1110011101000000",
    "1110011101011110",
    "1110101101101110",
    "1111001000111111",
    "1111100111000111",
    "1111111111100111",
    "1111101110000000",
    "1111100000100001",
    "1111010010100111",
    "1111000001100001",
    "1110101101000000",
    "1110011000010000",
    "1110001000011011",
    "1110000101000000",
    "1110010100101100",
    "1110110111011111",
    "1111100110101000",
    "1111101000101101",
    "1111000001110011",
    "1110101101010010",
    "1110110001100100",
    "1111001111001000",
    "1111111110100011",
    "1111001100000010",
    "1110011101001001",
    "1101111101111000",
    "1101110001111011",
    "1101110111110001",
    "1110001001001011",
    "1110011101110111",
    "1110101111001100",
    "1110111001111100",
    "1110111111000000",
    "1111000001111001",
    "1111000110001101",
    "1111001110101001",
    "1111011100101101",
    "1111110000011110",
    "1111110111100100",
    "1111011111010010",
    "1111001011101010",
    "1111000000011100",
    "1110111110111000",
    "1111000110100010",
    "1111010110000000",
    "1111101011000001",
    "1111111101000000",
    "1111100100110001",
    "1111001110001101",
    "1110111010100110",
    "1110101011010110",
    "1110100010000101",
    "1110100000001010",
    "1110100110100000",
    "1110110101001000",
    "1111001010111111",
    "1111100110000000",
    "1111111100110101",
    "1111100001010101",
    "1111001010110101",
    "1110111011100000",
    "1110110011111000",
    "1110110011001111",
    "1110111000100011",
    "1111000011000011",
    "1111010001111001",
    "1111100011101010",
    "1111110110000100",
    "1111111001110111",
    "1111101111001110",
    "1111101100100010",
    "1111110011100001",
    "1111111100000100",
    "1111100101011111",
    "1111001101100100",
    "1110111000111111",
    "1110101010100101",
    "1110100010110011",
    "1110100000001101",
    "1110100000000111",
    "1110011111111011",
    "1110011110111010",
    "1110011110000101",
    "1110011111101001",
    "1110100101100000",
    "1110101111110110",
    "1110111110101110",
    "1111010011100110",
    "1111101111001100",
    "1111101111100011",
    "1111001100001010",
    "1110101100001001",
    "1110010100111001",
    "1110001010100011",
    "1110001110101001",
    "1110011110000100",
    "1110110010010000",
    "1111000100100010",
    "1111001111011110",
    "1111010001010111",
    "1111001011111010",
    "1111000010100100",
    "1110111100001110",
    "1111000000011111",
    "1111010010100111",
    "1111110001000110",
    "1111101010010001",
    "1111001000011010",
    "1110110000000101",
    "1110100101000110",
    "1110100111001001",
    "1110110001100010",
    "1110111110110001",
    "1111001010001100",
    "1111010001000101",
    "1111010100000001",
    "1111010101110110",
    "1111011011000110",
    "1111100111110001",
    "1111111100000101",
    "1111101011011101",
    "1111010100011101",
    "1111000100011010",
    "1110111110110101",
    "1111000100001101",
    "1111010010001101",
    "1111100101000101",
    "1111111001101001",
    "1111110010010010",
    "1111100000100100",
    "1111010010101100",
    "1111001010000001",
    "1111000111001001",
    "1111001001101010",
    "1111010000010111",
    "1111011001001011",
    "1111100010101011",
    "1111101110100000",
    "1111111111000110",
    "1111101010011110",
    "1111001111000111",
    "1110110010011100",
    "1110011001101111",
    "1110001010001110",
    "1110000111111110",
    "1110010010100100",
    "1110100101100000",
    "1110111101001110",
    "1111011000100101",
    "1111110111110010",
    "1111100101001110",
    "1111000001010101",
    "1110100001101100",
    "1110001011101011",
    "1110000100001110",
    "1110001100110101",
    "1110100001010111",
    "1110111010111010",
    "1111010010011111",
    "1111100011000110",
    "1111101100100111",
    "1111110010111100",
    "1111111011010111",
    "1111110101110111",
    "1111100000100011",
    "1111001000010001",
    "1110110001110100",
    "1110100001111000",
    "1110011011010100",
    "1110011101111010",
    "1110100111001000",
    "1110110011011101",
    "1110111111111101",
    "1111001011001001",
    "1111010100001011",
    "1111011010001100",
    "1111011111000000",
    "1111100110111101",
    "1111110101011001",
    "1111110100110111",
    "1111011010011101",
    "1111000000100111",
    "1110101100101101",
    "1110100011000101",
    "1110100101011111",
    "1110110001001000",
    "1111000000100110",
    "1111001110011110",
    "1111010111100000",
    "1111011011100110",
    "1111011100010100",
    "1111011011010100",
    "1111011010000111",
    "1111011000110010",
    "1111010110011010",
    "1111010010011111",
    "1111001101011100",
    "1111001000110000",
    "1111000110100100",
    "1111001000011011",
    "1111001110010110",
    "1111010110100101",
    "1111011110101011",
    "1111100100110111",
    "1111101000101010",
    "1111101010001010",
    "1111101010000011",
    "1111101001100101",
    "1111101010001010",
    "1111101101100010",
    "1111110101110111",
    "1111111011101000",
    "1111100111011011",
    "1111001111110000",
    "1110111000100111",
    "1110100110110110",
    "1110011110010010",
    "1110100000010001",
    "1110101010110000",
    "1110111001010011",
    "1111000111011000",
    "1111010001010111",
    "1111010110011010",
    "1111011010011000",
    "1111100010111110",
    "1111110100000001",
    "1111110010111011",
    "1111010111010110",
    "1111000000111011",
    "1110110101111011",
    "1110111001100011",
    "1111001001110010",
    "1111011111110001",
    "1111110100000100",
    "1111111110101111",
    "1111111010100001",
    "1111111101000111",
    "1111111100110111",
    "1111111001000110",
    "1111111101111100",
    "1111110010001101",
    "1111011001011000",
    "1110111101000010",
    "1110100100101111",
    "1110010110010000",
    "1110010100001110",
    "1110011101100110",
    "1110101101001010",
    "1110111101000100",
    "1111001000011000",
    "1111001100010100",
    "1111001011110011",
    "1111001110000010",
    "1111011001001011",
    "1111110000010110",
    "1111101110110110",
    "1111001011110011",
    "1110101110010100",
    "1110011100111000",
    "1110011010001001",
    "1110100010100010",
    "1110101111110011",
    "1110111100001010",
    "1111000100011111",
    "1111001001001001",
    "1111001011110111",
    "1111001110011100",
    "1111010010111110",
    "1111011010000001",
    "1111100100011101",
    "1111110100100110",
    "1111110100111110",
    "1111011001100011",
    "1110111100001010",
    "1110100001111101",
    "1110001111111010",
    "1110001010001011",
    "1110010001100010",
    "1110100001011110",
    "1110110011010111",
    "1111000001000000",
    "1111001000010001",
    "1111001101010111",
    "1111010110010110",
    "1111100111000011",
    "1111111111101010",
    "1111100100110011",
    "1111001101111000",
    "1111000001110100",
    "1111000011110110",
    "1111010001000000",
    "1111100010000011",
    "1111110000000000",
    "1111110110011100",
    "1111110101000101",
    "1111101110111001",
    "1111100111000101",
    "1111100000000111",
    "1111011010101010",
    "1111010101011111",
    "1111010000110011",
    "1111001111001010",
    "1111010011011000",
    "1111011111011110",
    "1111110011000000",
    "1111110101110101",
    "1111100000101100",
    "1111010010101011",
    "1111001101111101",
    "1111010000011111",
    "1111010101101010",
    "1111011000110000",
    "1111010110001110",
    "1111001101110101",
    "1111000010000010",
    "1110110110000001",
    "1110101100110101",
    "1110101000000011",
    "1110101000011000",
    "1110101111000111",
    "1110111100101110",
    "1111010000010111",
    "1111100111101100",
    "1111111110110101",
    "1111101110100110",
    "1111100011111011",
    "1111100001110000",
    "1111100101001101",
    "1111101000110101",
    "1111100111001000",
    "1111011100111000",
    "1111001010111111",
    "1110110101110010",
    "1110100010110011",
    "1110010110100101",
    "1110010011000001",
    "1110010110111110",
    "1110011111011110",
    "1110101001001011",
    "1110110010101011",
    "1110111110001101",
    "1111001111100011",
    "1111101000110110",
    "1111110111000011",
    "1111010101001000",
    "1110110111101101",
    "1110100100001101",
    "1110011101010100",
    "1110100001101001",
    "1110101100011011",
    "1110110111111100",
    "1111000000110110",
    "1111001000100101",
    "1111010010110100",
    "1111100010010101",
    "1111110111101101",
    "1111101111100010",
    "1111011000000011",
    "1111000110111110",
    "1111000000110110",
    "1111000111010101",
    "1111011000101101",
    "1111110001001100",
    "1111110011111111",
    "1111011010111100",
    "1111000110100010",
    "1110111001000111",
    "1110110011011101",
    "1110110100100111",
    "1110111010011101",
    "1111000010100100",
    "1111001010110111",
    "1111010010101001",
    "1111011100100000",
    "1111101100101110",
    "1111111001101110",
    "1111010111000110",
    "1110110000011010",
    "1110001110010100",
    "1101111001000110",
    "1101110110010010",
    "1110000101010111",
    "1110011111101001",
    "1110111100001100",
    "1111010010111011",
    "1111011111001000",
    "1111100000111110",
    "1111011011001111",
    "1111010011111011",
    "1111010011000110",
    "1111011101100000",
    "1111110010101111",
    "1111110001110100",
    "1111011000010000",
    "1111000111011111",
    "1111000011011010",
    "1111001100010100",
    "1111011101110101",
    "1111110001010111",
    "1111111101000101",
    "1111101101001100",
    "1111011100000111",
    "1111000111101000",
    "1110110000101110",
    "1110011011000110",
    "1110001101011011",
    "1110010000101011",
    "1110101010000100",
    "1111010110110010",
    "1111110010111000",
    "1111000000011001",
    "1110011101000100",
    "1110001110001101",
    "1110010010100001",
    "1110100010100001",
    "1110110101001110",
    "1111000111001000",
    "1111011001011101",
    "1111101110111110",
    "1111110110010110",
    "1111011001000100",
    "1110111110011011",
    "1110101100011001",
    "1110101000000011",
    "1110110000110110",
    "1111000001001000",
    "1111010001111101",
    "1111011101011001",
    "1111100011000001",
    "1111101000001010",
    "1111110010111001",
    "1111111001000010",
    "1111011100110011",
    "1110111111000000",
    "1110100111101010",
    "1110011101000000",
    "1110100001010000",
    "1110110000101100",
    "1111000100111011",
    "1111011000010000",
    "1111100111000100",
    "1111110001000011",
    "1111110111001100",
    "1111111001110110",
    "1111111011000000",
    "1111111110100101",
    "1111111000001111",
    "1111101000000010",
    "1111010010010100",
    "1110111011101111",
    "1110101001011110",
    "1110100000010001",
    "1110100010110110",
    "1110101111010110",
    "1111000000011001",
    "1111001111100110",
    "1111010111100111",
    "1111010110110111",
    "1111001110110101",
    "1111000010111001",
    "1110110111101101",
    "1110110000010100",
    "1110101100110011",
    "1110101011110111",
    "1110101011101010",
    "1110101100101010",
    "1110110010001010",
    "1110111111010010",
    "1111010100111001",
    "1111110000011011",
    "1111110011000101",
    "1111011010101000",
    "1111001001011001",
    "1111000000000000",
    "1110111100001001",
    "1110111010011110",
    "1110111000100010",
    "1110110101100100",
    "1110110010110011",
    "1110110001111011",
    "1110110100000110",
    "1110111010100101",
    "1111000110100100",
    "1111011000010001",
    "1111101110101011",
    "1111111001001110",
    "1111100011100110",
    "1111010011110110",
    "1111001100011100",
    "1111001110100011",
    "1111011001010001",
    "1111101001111110",
    "1111111101000000",
    "1111110001011000",
    "1111100011101110",
    "1111011010111111",
    "1111010111011010",
    "1111011000100000",
    "1111011110001101",
    "1111101000100001",
    "1111110111000111",
    "1111110110101000",
    "1111100010011100",
    "1111001111000010",
    "1110111111110001",
    "1110110111101010",
    "1110110111101010",
    "1110111110011001",
    "1111001001010000",
    "1111010100110110",
    "1111011110010001",
    "1111100011101001",
    "1111100100111011",
    "1111100011110100",
    "1111100010110100",
    "1111100101001110",
    "1111101111000101",
    "1111111101101001",
    "1111100010000110",
    "1111000010100001",
    "1110100101001001",
    "1110010000001100",
    "1110001000000100",
    "1110001110001101",
    "1110100001100100",
    "1111000000110110",
    "1111101001010010",
    "1111101001111101",
    "1110111110111010",
    "1110011100010100",
    "1110000111101100",
    "1110000011100111",
    "1110001111100100",
    "1110100110011111",
    "1111000000011110",
    "1111010110011011",
    "1111100011100111",
    "1111100111110100",
    "1111101000110111",
    "1111101110110000",
    "1111111111101100",
    "1111100011000000",
    "1110111110101011",
    "1110011011110111",
    "1110000010110110",
    "1101111001010001",
    "1101111110011011",
    "1110001100011110",
    "1110011100101110",
    "1110101010100010",
    "1110110110110010",
    "1111000110010110",
    "1111011100100001",
    "1111111001101011",
    "1111100110000011",
    "1111001010011001",
    "1110111010010110",
    "1110111010000100",
    "1111001000101010",
    "1111011111001101",
    "1111110101000100",
    "1111111100100101",
    "1111111000100100",
    "1111111011111000",
    "1111111111110011",
    "1111111110000000",
    "1111110010111100",
    "1111011111011110",
    "1111001000011101",
    "1110110011100001",
    "1110100101011101",
    "1110100001010100",
    "1110100110000000",
    "1110101111110001",
    "1110111100101101",
    "1111001101110011",
    "1111100100100100",
    "1111111111000100",
    "1111100000011111",
    "1111000100111100",
    "1110110001101110",
    "1110101011100001",
    "1110110011011000",
    "1111000101101110",
    "1111011100101011",
    "1111110010111000",
    "1111111001011101",
    "1111100110110101",
    "1111010011011010",
    "1110111110100110",
    "1110101010000010",
    "1110011001011101",
    "1110010000110001",
    "1110010010010100",
    "1110011101010001",
    "1110101101011001",
    "1110111101101000",
    "1111001001111111",
    "1111010001011010",
    "1111010101100101",
    "1111011001001001",
    "1111011111011001",
    "1111101011100000",
    "1111111110001001",
    "1111101010101111",
    "1111010011011010",
    "1111000000101100",
    "1110110110010101",
    "1110110110001000",
    "1111000000010101",
    "1111010100011000",
    "1111110000100100",
    "1111101101101100",
    "1111001010000111",
    "1110101001010101",
    "1110010000000101",
    "1110000010001011",
    "1110000001001000",
    "1110001011001001",
    "1110011011111010",
    "1110101110111010",
    "1111000001111110",
    "1111010101100111",
    "1111101011000110",
    "1111111101010001",
    "1111100100110011",
    "1111001110000100",
    "1110111100001100",
    "1110110001111000",
    "1110101111110011",
    "1110110100010101",
    "1110111100010110",
    "1111000100100000",
    "1111001011000010",
    "1111010000001100",
    "1111010101011111",
    "1111011100100011",
    "1111100101110010",
    "1111101111011000",
    "1111110101101000",
    "1111110100101100",
    "1111101010010110",
    "1111010111010001",
    "1110111111011010",
    "1110101000101010",
    "1110011000010001",
    "1110010001010101",
    "1110010100001110",
    "1110011111000101",
    "1110101110101000",
    "1110111111010001",
    "1111001110011111",
    "1111011011010110",
    "1111100110001000",
    "1111101111100100",
    "1111111000010101",
    "1111111110111110",
    "1111110110010111",
    "1111101110111010",
    "1111101010110011",
    "1111101100010111",
    "1111110101000101",
    "1111111011011100",
    "1111100111100011",
    "1111010010101110",
    "1111000000101110",
    "1110110100011100",
    "1110101110110000",
    "1110101110101011",
    "1110110011100111",
    "1110111110110110",
    "1111010010010100",
    "1111101110011100",
    "1111101111001101",
    "1111001100001001",
    "1110101110110110",
    "1110011100101011",
    "1110011000001000",
    "1110011110111111",
    "1110101100101010",
    "1110111110101110",
    "1111010101000000",
    "1111110000000110",
    "1111101111111011",
    "1111001110000100",
    "1110101111001111",
    "1110011001001011",
    "1110010001001010",
    "1110011000001110",
    "1110101010100101",
    "1111000100100100",
    "1111100100000000",
    "1111111000100100",
    "1111010010000110",
    "1110101011000111",
    "1110000111110101",
    "1101101100100011",
    "1101011101110010",
    "1101011101101011",
    "1101101001101101",
    "1101111101000010",
    "1110010010010100",
    "1110100101001001",
    "1110110100001010",
    "1111000001001111",
    "1111010001110110",
    "1111101011010111",
    "1111110001010000",
    "1111001000101100",
    "1110100011000101",
    "1110001001010000",
    "1110000001001100",
    "1110001100000111",
    "1110100100111011",
    "1111000010101011",
    "1111011101000111",
    "1111101110111011",
    "1111110110111110",
    "1111110111011001",
    "1111110011100101",
    "1111101110111010",
    "1111101011011001",
    "1111101000101100",
    "1111100101101010",
    "1111100001101001",
    "1111011100100110",
    "1111010111100111",
    "1111010011111011",
    "1111010011010010",
    "1111011000100011",
    "1111100110011000",
    "1111111101100001",
    "1111100011010011",
    "1111000000100111",
    "1110100000100100",
    "1110001000111010",
    "1101111101010110",
    "1101111101000111",
    "1110000011111000",
    "1110001100101110",
    "1110010011101100",
    "1110010111100101",
    "1110011100010001",
    "1110100111111001",
    "1110111110101000",
    "1111100000101110",
    "1111110110111001",
    "1111010000011010",
    "1110110011010011",
    "1110100101001110",
    "1110100110100111",
    "1110110010000110",
    "1111000000100100",
    "1111001011111101",
    "1111010001000011",
    "1111010000010101",
    "1111001011110011",
    "1111000110000000",
    "1111000001011010",
    "1110111110110101",
    "1110111111101001",
    "1111000110011101",
    "1111010100101010",
    "1111101010000110",
    "1111111011000111",
    "1111011110110110",
    "1111000101100111",
    "1110110011110001",
    "1110101011011001",
    "1110101010100110",
    "1110101101100001",
    "1110110000010101",
    "1110110000100011",
    "1110101110000010",
    "1110101010001110",
    "1110100110101010",
    "1110100101010010",
    "1110101000101100",
    "1110110011100010",
    "1111000111000110",
    "1111100010011010",
    "1111111101110111",
    "1111011110110001",
    "1111000101100101",
    "1110111000001100",
    "1110111010101010",
    "1111001100011001",
    "1111101000111110",
    "1111110110101000",
    "1111011010001100",
    "1111000110111001",
    "1110111111000111",
    "1111000001110011",
    "1111001010100010",
    "1111010100101010",
    "1111011100110011",
    "1111100010100111",
    "1111101010011001",
    "1111111000101001",
    "1111110001010110",
    "1111010110000110",
    "1110111011101111",
    "1110101001010101",
    "1110100100000011",
    "1110101101110011",
    "1111000010100110",
    "1111011010111000",
    "1111110010001010",
    "1111111000010010",
    "1111100010110110",
    "1111001011011011",
    "1110110010110001",
    "1110011100000010",
    "1110001011011000",
    "1110000101010000",
    "1110001011010100",
    "1110011011010001",
    "1110110000111101",
    "1111001001001100",
    "1111100100000001",
    "1111111100100000",
    "1111010111101111",
    "1110101111101011",
    "1110001001100011",
    "1101101100100000",
    "1101011110011110",
    "1101100001111000",
    "1101110011111000",
    "1110001101100110",
    "1110100111001011",
    "1110111010010001",
    "1111000100011000",
    "1111000110100100",
    "1111000011001101",
    "1110111101010010",
    "1110110110110010",
    "1110110000100001",
    "1110101101000101",
    "1110110000111000",
    "1110111110110001",
    "1111010111001000",
    "1111110110110001",
    "1111101000100111",
    "1111001110011100",
    "1111000000110011",
    "1111000001111011",
    "1111001101101001",
    "1111011100101010",
    "1111101000001010",
    "1111101011011100",
    "1111100111000100",
    "1111100001101001",
    "1111100011000000",
    "1111110000100111",
    "1111110101011001",
    "1111010101010010",
    "1110110111011101",
    "1110100011010000",
    "1110011100110011",
    "1110100001111110",
    "1110101101100001",
    "1110111011111000",
    "1111001011101111",
    "1111011101100011",
    "1111110001101000",
    "1111111010011111",
    "1111101010100011",
    "1111100010111011",
    "1111100111011110",
    "1111110111110001",
    "1111110000101100",
    "1111011000011101",
    "1111000110001101",
    "1110111101101101",
    "1110111110111010",
    "1111000110101101",
    "1111010000001100",
    "1111010111010011",
    "1111011010110101",
    "1111011100101110",
    "1111100010010000",
    "1111110000101000",
    "1111110110101110",
    "1111010110101101",
    "1110110101011000",
    "1110011001110101",
    "1110001001100010",
    "1110000111001001",
    "1110010001000000",
    "1110100010000011",
    "1110110100110100",
    "1111000100111011",
    "1111010000011100",
    "1111010111111111",
    "1111011100111111",
    "1111100000110001",
    "1111100101001101",
    "1111101100110001",
    "1111111001101010",
    "1111110011101010",
    "1111011101111000",
    "1111001001010110",
    "1110111010101011",
    "1110110101001000",
    "1110111001100011",
    "1111000101100100",
    "1111010011111110",
    "1111011111010100",
    "1111100100000110",
    "1111100010000000",
    "1111011011001111",
    "1111010011001101",
    "1111001100111000",
    "1111001001110100",
    "1111001001101111",
    "1111001011100000",
    "1111001101110010",
    "1111001111110011",
    "1111010011011000",
    "1111011101000010",
    "1111110000000111",
    "1111110011101010",
    "1111010010110011",
    "1110110100011000",
    "1110011111001000",
    "1110010111110111",
    "1110011111101000",
    "1110110010001111",
    "1111001000011000",
    "1111011011111100",
    "1111101100000001",
    "1111111100011111",
    "1111101110100100",
    "1111010100001011",
    "1110110111100000",
    "1110011110111101",
    "1110010001001000",
    "1110010010101100",
    "1110100011001010",
    "1110111100100011",
    "1111011000111111",
    "1111110101111111",
    "1111101100100011",
    "1111001101100001",
    "1110101101111000",
    "1110010001011001",
    "1101111100010110",
    "1101110011000110",
    "1101110111100010",
    "1110000110011000",
    "1110011011111101",
    "1110110110100101",
    "1111010100110110",
    "1111110101101101",
    "1111101000111101",
    "1111001011011011",
    "1110110101111001",
    "1110101100111010",
    "1110110011000011",
    "1111000100111001",
    "1111011011110011",
    "1111110000111001",
    "1111111110101101",
    "1111111010101011",
    "1111110110110100",
    "1111110000111000",
    "1111100101101001",
    "1111010110011000",
    "1111001000100111",
    "1111000001111110",
    "1111000111000011",
    "1111011001010110",
    "1111110101010100",
    "1111101010101001",
    "1111001011101011",
    "1110110001011010",
    "1110011101100000",
    "1110010000101001",
    "1110001011001100",
    "1110001100010110",
    "1110010011100010",
    "1110100000100011",
    "1110110001111101",
    "1111000101110100",
    "1111011001011000",
    "1111101010001011",
    "1111111010001000",
    "1111110010100001",
    "1111011001000110",
    "1110111001101000",
    "1110011000110101",
    "1101111101111010",
    "1101101111000101",
    "1101110000001010",
    "1101111111011100",
    "1110010110000011",
    "1110101100010011",
    "1110111100011100",
    "1111000100000110",
    "1111000101000101",
    "1111000101001101",
    "1111001011110011",
    "1111011101001111",
    "1111111000010010",
    "1111101000110000",
    "1111001101100000",
    "1110111100001010",
    "1110110111101111",
    "1110111110000111",
    "1111001001000110",
    "1111010010110100",
    "1111011000000110",
    "1111011000001001",
    "1111010101000101",
    "1111010100001010",
    "1111011011100000",
    "1111101110100100",
    "1111110011110011",
    "1111010001011111",
    "1110110001111110",
    "1110011011101111",
    "1110010010100110",
    "1110010101110001",
    "1110100000111101",
    "1110110000100100",
    "1111000010101011",
    "1111010110001011",
    "1111101010000101",
    "1111111011100100",
    "1111111001000100",
    "1111110110111010",
    "1111111111101000",
    "1111101110011101",
    "1111011000111001",
    "1111000101111110",
    "1110111011011001",
    "1110111100001001",
    "1111000111001011",
    "1111011000101111",
    "1111101011011010",
    "1111111010011001",
    "1111111100001100",
    "1111110111010110",
    "1111110100110100",
    "1111110001110110",
    "1111101011110110",
    "1111100001000111",
    "1111010001010111",
    "1110111110011001",
    "1110101011011110",
    "1110011100000111",
    "1110010011000101",
    "1110010001111011",
    "1110011000010101",
    "1110100100001000",
    "1110110011011101",
    "1111000110100000",
    "1111011110000101",
    "1111111001101001",
    "1111101001001010",
    "1111001101111011",
    "1110111000011000",
    "1110101011110101",
    "1110101010010110",
    "1110110011110110",
    "1111000110101010",
    "1111100000001000",
    "1111111100110011",
    "1111100111000011",
    "1111001111010111",
    "1110111111101001",
    "1110111001100010",
    "1110111101101001",
    "1111001101000000",
    "1111100110101111",
    "1111111000011000",
    "1111010101010111",
    "1110110110011101",
    "1110100001001010",
    "1110011000100111",
    "1110011101000111",
    "1110101011001100",
    "1110111101001100",
    "1111001111110101",
    "1111100011101001",
    "1111111010110100",
    "1111101001001101",
    "1111001010000110",
    "1110101100010111",
    "1110010101001001",
    "1110001001011001",
    "1110001011100000",
    "1110011000110100",
    "1110101011110010",
    "1110111110111000",
    "1111001110000100",
    "1111011000100111",
    "1111100000001111",
    "1111100111000000",
    "1111101111000001",
    "1111111001101001",
    "1111111000111001",
    "1111101001011111",
    "1111011010001110",
    "1111001101111000",
    "1111000110011111",
    "1111000100111110",
    "1111001001010000",
    "1111010001111011",
    "1111011100100001",
    "1111100101110110",
    "1111101011001110",
    "1111101011110000",
    "1111101000000100",
    "1111100001100010",
    "1111011010000100",
    "1111010011010010",
    "1111001110001101",
    "1111001011000001",
    "1111001000111100",
    "1111000110110110",
    "1111000011111110",
    "1111000000000111",
    "1110111101011001",
    "1111000000111001",
    "1111001110110110",
    "1111101000010101",
    "1111110101110001",
    "1111010010111001",
    "1110110111000011",
    "1110101000010001",
    "1110101000011110",
    "1110110011011100",
    "1111000001100010",
    "1111001100010100",
    "1111010000010001",
    "1111001110001010",
    "1111001001101111",
    "1111000110010110",
    "1111000111010101",
    "1111010000100001",
    "1111100011100010",
    "1111111111000110",
    "1111100000010111",
    "1111000000111001",
    "1110101000010101",
    "1110011010110010",
    "1110011010010011",
    "1110100101000001",
    "1110110101101001",
    "1111000110100100",
    "1111010010111101",
    "1111011001100000",
    "1111011110110101",
    "1111101000111000",
    "1111111011100110",
    "1111101000101001",
    "1111001001010001",
    "1110101101100110",
    "1110011100001010",
    "1110011010110100",
    "1110101010111111",
    "1111001000010110",
    "1111101100001100",
    "1111110000110111",
    "1111010100101010",
    "1111000001111110",
    "1110111001111111",
    "1110111010111100",
    "1111000000011100",
    "1111000110110100",
    "1111001011110111",
    "1111001110111111",
    "1111010001011110",
    "1111010100011101",
    "1111011000100101",
    "1111011110100011",
    "1111100110010010",
    "1111101110101111",
    "1111110110010111",
    "1111111010110110",
    "1111111010011001",
    "1111110100111011",
    "1111101011011001",
    "1111011111101001",
    "1111010011110110",
    "1111001001111010",
    "1111000011010111",
    "1111000001000011",
    "1111000100100100",
    "1111010000001000",
    "1111100101010010",
    "1111111100100000",
    "1111011000011011",
    "1110110100000001",
    "1110010101010111",
    "1110000001011100",
    "1101111010101000",
    "1101111111010010",
    "1110001011000110",
    "1110011000101000",
    "1110100011011101",
    "1110101001110111",
    "1110101100100110",
    "1110101101011011",
    "1110101110000010",
    "1110110000110000",
    "1110111001010001",
    "1111001010001100",
    "1111100011001101",
    "1111111110111010",
    "1111100010000000",
    "1111001011100110",
    "1110111111110001",
    "1111000000000000",
    "1111001001011001",
    "1111010110111011",
    "1111100011011100",
    "1111101100100000",
    "1111110101010010",
    "1111111101001111",
    "1111101000111011",
    "1111001111001100",
    "1110110101101110",
    "1110100011100010",
    "1110011101111010",
    "1110100110101010",
    "1110111001111101",
    "1111001111101001",
    "1111011111110110",
    "1111100101100010",
    "1111100000110011",
    "1111010101011000",
    "1111000111011011",
    "1110111100010100",
    "1110111010000001",
    "1111000011100111",
    "1111011000100011",
    "1111110100110101",
    "1111101110001001",
    "1111010110101100",
    "1111001000111111",
    "1111000110100101",
    "1111001101011100",
    "1111011001001100",
    "1111100100111011",
    "1111101100101100",
    "1111110001011100",
    "1111110111111101",
    "1111111011110000",
    "1111101000000101",
    "1111001111001100",
    "1110110111001001",
    "1110100110010010",
    "1110100001010101",
    "1110101001010000",
    "1110111001000001",
    "1111001001010101",
    "1111010100000110",
    "1111010110011010",
    "1111010010000101",
    "1111001010110100",
    "1111000100001110",
    "1111000011010010",
    "1111001100010100",
    "1111011111111011",
    "1111111011010011",
    "1111100111101101",
    "1111010000000101",
    "1111000001111001",
    "1110111110101101",
    "1111000101000001",
    "1111010000000010",
    "1111011010011001",
    "1111100010001000",
    "1111101000111000",
    "1111110010001111",
    "1111111111010011",
    "1111101101001101",
    "1111011011001100",
    "1111001110001010",
    "1111001010110000",
    "1111010010000010",
    "1111100000100100",
    "1111110000111100",
    "1111111101001101",
    "1111111110101001",
    "1111111110111001",
    "1111111101000000",
    "1111111100101111",
    "1111101010011001",
    "1111001101101001",
    "1110101101010110",
    "1110010001111000",
    "1110000010110110",
    "1110000100010000",
    "1110010011100100",
    "1110101001101010",
    "1110111111001100",
    "1111001110101110",
    "1111010111010000",
    "1111011101001110",
    "1111100110010110",
    "1111110110110101",
    "1111110001000001",
    "1111010110011011",
    "1111000000011100",
    "1110110101010000",
    "1110111000001000",
    "1111000110100010",
    "1111011001011110",
    "1111101010000100",
    "1111110011100100",
    "1111110100110011",
    "1111101111110011",
    "1111100111011100",
    "1111011111000101",
    "1111011001101111",
    "1111011000001011",
    "1111011001110010",
    "1111011101001111",
    "1111100000011111",
    "1111100010100110",
    "1111100100001011",
    "1111100110110100",
    "1111101011010001",
    "1111110000100100",
    "1111110100010011",
    "1111110011111100",
    "1111101110001000",
    "1111100011010011",
    "1111010110001101",
    "1111001010011000",
    "1111000011000000",
    "1111000001111011",
    "1111000110111111",
    "1111010000001101",
    "1111011010101101",
    "1111100100100010",
    "1111101111000111",
    "1111111101111110",
    "1111101100001101",
    "1111001111011010",
    "1110101111001010",
    "1110010001010000",
    "1101111011001111",
    "1101110000111101",
    "1101110010011100",
    "1101111011110101",
    "1110001000011011",
    "1110010011110011",
    "1110011100011110",
    "1110100110010011",
    "1110110110001011",
    "1111001110110000",
    "1111101111010110",
    "1111101101100100",
    "1111001111100001",
    "1110111100110111",
    "1110111001100010",
    "1111000100010000",
    "1111010111011000",
    "1111101100110010",
    "1111111111100010",
    "1111110000111100",
    "1111100000111000",
    "1111001100101101",
    "1110110011000101",
    "1110010101101110",
    "1101111010010110",
    "1101100111000001",
    "1101100000001100",
    "1101100111011101",
    "1101111001010001",
    "1110001111011100",
    "1110100100001011",
    "1110110011101110",
    "1110111101010001",
    "1111000010011010",
    "1111000111010110",
    "1111010001011010",
    "1111100011100100",
    "1111111101000110",
    "1111100110000000",
    "1111001100000010",
    "1110111010111010",
    "1110110110100010",
    "1110111111000000",
    "1111010000010010",
    "1111100100110001",
    "1111110111011001",
    "1111111010011000",
    "1111110000010010",
    "1111101000111101",
    "1111100011011000",
    "1111011111010001",
    "1111011101010010",
    "1111011110010100",
    "1111100010011010",
    "1111101000001010",
    "1111101100101001",
    "1111101100011010",
    "1111100101101111",
    "1111011001110101",
    "1111001101000010",
    "1111000101101100",
    "1111001001000111",
    "1111011001000010",
    "1111110010111110",
    "1111101110101010",
    "1111010010101011",
    "1110111110110001",
    "1110110110101100",
    "1110111010010011",
    "1111000101111110",
    "1111010101001001",
    "1111100011111100",
    "1111101111101010",
    "1111110111101010",
    "1111111100111100",
    "1111111110110000",
    "1111111010100000",
    "1111110111011110",
    "1111111000001100",
    "1111111110101011",
    "1111110100000101",
    "1111100001010111",
    "1111001100100000",
    "1110111001110010",
    "1110101100111000",
    "1110100111011010",
    "1110101000101101",
    "1110101110001101",
    "1110110101010101",
    "1110111101111011",
    "1111001010000010",
    "1111011011110011",
    "1111110011111101",
    "1111101111001100",
    "1111010001011010",
    "1110110111010001",
    "1110100101000110",
    "1110011100100011",
    "1110011011110101",
    "1110011111011111",
    "1110100011111011",
    "1110100111000100",
    "1110101000101111",
    "1110101001011101",
    "1110101100100000",
    "1110110110111111",
    "1111001011101111",
    "1111101010000101",
    "1111110010100010",
    "1111010001100110",
    "1110111001101010",
    "1110101110111000",
    "1110110001010111",
    "1110111101111101",
    "1111010001110000",
    "1111101001011110",
    "1111111110010010",
    "1111101000000101",
    "1111010110100100",
    "1111001100000001",
    "1111001011000001",
    "1111010110111110",
    "1111110000001111",
    "1111101100110011",
    "1111000110011111",
    "1110100100101110",
    "1110001110000010",
    "1110000110010011",
    "1110001101100001",
    "1110011110111000",
    "1110110011100010",
    "1111000110011101",
    "1111010111001011",
    "1111101001000110",
    "1111111111011011",
    "1111100101000110",
    "1111000110111110",
    "1110101011000111",
    "1110010110011011",
    "1110001100110000",
    "1110001110111010",
    "1110011001101011",
    "1110101000000100",
    "1110110110000011",
    "1111000011010000",
    "1111010010010101",
    "1111100100111100",
    "1111111001101011",
    "1111110011101110",
    "1111101001001000",
    "1111101010100111",
    "1111111000000111",
    "1111110011111001",
    "1111100010001011",
    "1111011010101011",
    "1111100001100111",
    "1111110100110110",
    "1111110010010111",
    "1111011011001010",
    "1111001010100000",
    "1111000001101100",
    "1110111110100001",
    "1110111101101000",
    "1110111100000100",
    "1110111001010000",
    "1110110111101101",
    "1110111010111100",
    "1111000100101001",
    "1111010010111001",
    "1111100000100111",
    "1111101000100110",
    "1111101000000101",
    "1111011111011111",
    "1111010010101001",
    "1111000111011101",
    "1111000011101110",
    "1111001011000111",
    "1111011101101000",
    "1111110111010101",
    "1111101101110100",
    "1111010111100111",
    "1111001010001100",
    "1111000111011011",
    "1111001110111011",
    "1111011110001101",
    "1111110001011000",
    "1111111011100100",
    "1111101100000001",
    "1111100010100100",
    "1111100001000111",
    "1111101000001110",
    "1111110110011111",
    "1111110111101000",
    "1111100110100101",
    "1111011010000110",
    "1111010100011101",
    "1111010101111011",
    "1111011101000101",
    "1111100111101010",
    "1111110010101000",
    "1111111011010000",
    "1111111111101001",
    "1111111111001101",
    "1111111010101000",
    "1111110011011000",
    "1111101011100111",
    "1111100101101111",
    "1111100100010111",
    "1111101001101111",
    "1111110110100001",
    "1111110110111000",
    "1111100010000101",
    "1111001111011001",
    "1111000010101111",
    "1110111110000101",
    "1111000001110110",
    "1111001110010100",
    "1111100010110100",
    "1111111100111101",
    "1111100111001000",
    "1111001110100100",
    "1110111101111011",
    "1110110111110101",
    "1110111100100000",
    "1111001000100101",
    "1111010110100111",
    "1111100001110000",
    "1111100110110101",
    "1111100101010011",
    "1111100000001111",
    "1111011110000111",
    "1111100101100111",
    "1111111010000101",
    "1111100110001101",
    "1111000001111101",
    "1110100001010010",
    "1110001011001010",
    "1110000011010011",
    "1110001000000110",
    "1110010100101001",
    "1110100100000011",
    "1110110010110110",
    "1110111111101100",
    "1111001010011101",
    "1111010100100111",
    "1111100010000110",
    "1111110101100011",
    "1111110001011111",
    "1111010110100000",
    "1110111111001101",
    "1110110000111101",
    "1110101110110001",
    "1110111000011101",
    "1111001001100011",
    "1111011100001110",
    "1111101011001101",
    "1111110100110101",
    "1111111100110011",
    "1111110111101111",
    "1111100101100111",
    "1111001100010110",
    "1110110000000000",
    "1110010111001101",
    "1110001000010000",
    "1110001001000100",
    "1110011100000111",
    "1110111110010111",
    "1111101001011011",
    "1111101011001100",
    "1111000111001011",
    "1110101111001000",
    "1110100101111001",
    "1110101010110101",
    "1110111000110100",
    "1111001011011101",
    "1111100001110110",
    "1111111100001010",
    "1111100101000110",
    "1111000100001000",
    "1110100110011010",
    "1110010001000111",
    "1110001000010110",
    "1110001101101110",
    "1110011111001111",
    "1110111010101010",
    "1111011100110011",
    "1111111110101111",
    "1111011011110111",
    "1110111110011001",
    "1110101001001100",
    "1110011101000100",
    "1110011010001110",
    "1110011111011010",
    "1110101011001010",
    "1110111101101001",
    "1111010110011010",
    "1111110011100110",
    "1111101101100111",
    "1111010001011001",
    "1110111010100110",
    "1110101011001100",
    "1110100100010010",
    "1110100100101111",
    "1110101001111010",
    "1110110000110001",
    "1110110110101101",
    "1110111010110000",
    "1110111101011100",
    "1111000001001101",
    "1111001010000001",
    "1111011010100110",
    "1111110010101100",
    "1111110000100010",
    "1111010011111100",
    "1110111101010001",
    "1110110000110101",
    "1110110000011001",
    "1110111010010110",
    "1111001010001001",
    "1111011010011001",
    "1111100110101111",
    "1111101100100111",
    "1111101011111100",
    "1111100110011010",
    "1111011110011111",
    "1111010111001110",
    "1111010011001000",
    "1111010100001110",
    "1111011011100110",
    "1111101000011000",
    "1111111000010001",
    "1111110111011000",
    "1111101001000001",
    "1111011110000100",
    "1111010111011101",
    "1111010110001000",
    "1111011010101000",
    "1111100100110100",
    "1111110011000011",
    "1111111110000001",
    "1111110010010101",
    "1111101100111100",
    "1111101111010111",
    "1111111000111000",
    "1111111000111001",
    "1111101001010110",
    "1111011011100101",
    "1111010001101001",
    "1111001100000001",
    "1111001010000010",
    "1111001010010001",
    "1111001011001010",
    "1111001011110101",
    "1111001100000101",
    "1111001011111010",
    "1111001011010110",
    "1111001010011011",
    "1111001001011101",
    "1111001001010110",
    "1111001011000100",
    "1111001111011110",
    "1111010110100100",
    "1111011111011111",
    "1111101000110101",
    "1111110000111110",
    "1111111000100101",
    "1111111101011110",
    "1111101111000110",
    "1111011100001001",
    "1111000111010000",
    "1110110101011010",
    "1110101011011001",
    "1110101100001111",
    "1110110111110001",
    "1111001001010101",
    "1111011011011011",
    "1111101011100001",
    "1111111001111010",
    "1111110111010000",
    "1111100110010011",
    "1111010100001011",
    "1111000011100010",
    "1110111000010000",
    "1110110110001000",
    "1110111101000101",
    "1111001001101010",
    "1111010111010110",
    "1111100001101110",
    "1111100110110010",
    "1111100111101010",
    "1111100110100001",
    "1111100110001110",
    "1111101000010001",
    "1111101100110011",
    "1111110101111100",
    "1111111010000101",
    "1111100011010011",
    "1111000111100000",
    "1110101011001100",
    "1110010011111011",
    "1110000110101100",
    "1110000110110100",
    "1110010010110011",
    "1110100100110001",
    "1110110110001001",
    "1111000001110000",
    "1111000101100101",
    "1111000101100000",
    "1111001000110010",
    "1111010101011111",
    "1111101110000011",
    "1111110001010110",
    "1111010000111101",
    "1110111000110101",
    "1110101111000000",
    "1110110100001011",
    "1111000010110110",
    "1111010011011101",
    "1111100000000011",
    "1111100101111011",
    "1111100110010011",
    "1111100100000110",
    "1111100001111001",
    "1111100001111101",
    "1111100100010111",
    "1111101000101111",
    "1111101111101111",
    "1111111010001100",
    "1111110111010011",
    "1111100100110011",
    "1111001111100011",
    "1110111010001011",
    "1110100111111100",
    "1110011011100000",
    "1110010101010010",
    "1110010011101001",
    "1110010100010101",
    "1110010101101001",
    "1110010111000001",
    "1110011000110111",
    "1110011011011110",
    "1110011110111101",
    "1110100011001111",
    "1110101000001000",
    "1110101101110101",
    "1110110100110011",
    "1110111100111000",
    "1111000101000110",
    "1111001011110011",
    "1111001111101000",
    "1111010000010100",
    "1111001111010111",
    "1111010000000011",
    "1111010110101000",
    "1111100101101010",
    "1111111100111110",
    "1111100110010000",
    "1111001001000001",
    "1110110000100100",
    "1110100000111011",
    "1110011011100110",
    "1110011111001101",
    "1110101000011000",
    "1110110011011010",
    "1110111101110010",
    "1111000110010110",
    "1111001101001010",
    "1111010011001101",
    "1111011001100011",
    "1111100000100110",
    "1111101001111110",
    "1111111000100101",
    "1111110010000110",
    "1111010110111110",
    "1110111001110111",
    "1110100000101011",
    "1110010000111000",
    "1110001110001101",
    "1110011000101010",
    "1110101011101000",
    "1111000001000101",
    "1111010011100111",
    "1111100000100100",
    "1111101010000101",
    "1111110100100111",
    "1111111100011001",
    "1111101000100100",
    "1111010011101110",
    "1111000100010011",
    "1110111111110001",
    "1111001000111001",
    "1111011101100000",
    "1111110110010111",
    "1111110101000101",
    "1111101011011011",
    "1111101110110001",
    "1111111100101011",
    "1111101111100111",
    "1111011011101011",
    "1111001100111111",
    "1111000111000011",
    "1111001010101011",
    "1111010110001110",
    "1111100110001101",
    "1111110110110001",
    "1111111010110010",
    "1111110000010001",
    "1111101010010010",
    "1111101000100110",
    "1111101010010101",
    "1111101110000000",
    "1111110001110101",
    "1111110100001101",
    "1111110011101111",
    "1111101111110001",
    "1111101000101011",
    "1111011111100100",
    "1111010110000100",
    "1111001101101011",
    "1111000111100000",
    "1111000100100111",
    "1111000101101100",
    "1111001011111100",
    "1111011001111001",
    "1111110000111011",
    "1111110000010010",
    "1111001110000111",
    "1110101111010010",
    "1110011010011000",
    "1110010011011000",
    "1110011010101000",
    "1110101011001001",
    "1110111101100011",
    "1111001101111011",
    "1111011100110111",
    "1111101101001101",
    "1111111110010101",
    "1111100110010110",
    "1111001110010001",
    "1110111010110100",
    "1110110001010000",
    "1110110100000000",
    "1111000010001101",
    "1111011001000111",
    "1111110011001101",
    "1111110110101110",
    "1111101011001000",
    "1111101101110001",
    "1111111110000000",
    "1111101000111011",
    "1111001101111111",
    "1110111000010110",
    "1110101110100001",
    "1110110100100111",
    "1111001010100010",
    "1111101011111010",
    "1111101101111001",
    "1111001010100110",
    "1110110000100100",
    "1110100010111001",
    "1110100000110101",
    "1110100101110100",
    "1110101100001001",
    "1110110000110001",
    "1110110101010101",
    "1110111101111101",
    "1111001101110000",
    "1111100100101110",
    "1111111111110100",
    "1111100101101100",
    "1111010001001000",
    "1111000110001011",
    "1111000100011101",
    "1111001001000010",
    "1111010010000110",
    "1111011111000100",
    "1111110000000101",
    "1111111010101000",
    "1111100011011000",
    "1111001110110001",
    "1111000010101110",
    "1111000100110111",
    "1111010110110110",
    "1111110100111111",
    "1111100111010000",
    "1111000110000100",
    "1110101110000101",
    "1110100010001101",
    "1110100001110100",
    "1110101001100101",
    "1110110101011000",
    "1111000010000011",
    "1111001101100110",
    "1111010111001110",
    "1111011111011111",
    "1111100111001000",
    "1111101110110001",
    "1111111001000110",
    "1111110110011000",
    "1111011110010001",
    "1110111111111111",
    "1110100000111001",
    "1110000111111110",
    "1101111010101000",
    "1101111011110010",
    "1110001001101011",
    "1110011110011011",
    "1110110011101111",
    "1111000101001001",
    "1111010001100100",
    "1111011011110011",
    "1111100111011010",
    "1111110111001110",
    "1111110100011010",
    "1111011111000111",
    "1111001110001010",
    "1111000110010011",
    "1111001001001011",
    "1111010100001000",
    "1111100001111011",
    "1111101101011001",
    "1111110011100000",
    "1111110100011000",
    "1111110001111111",
    "1111101110111001",
    "1111101100100110",
    "1111101100001011",
    "1111110000001011",
    "1111111011010000",
    "1111110001110010",
    "1111011000100101",
    "1110111101100000",
    "1110100101101110",
    "1110010101111001",
    "1110010001000010",
    "1110010110000000",
    "1110100000010001",
    "1110101010100010",
    "1110110000100011",
    "1110110000110101",
    "1110101100110000",
    "1110100111101101",
    "1110100110100010",
    "1110101110000111",
    "1111000000100110",
    "1111011101000000",
    "1111111111100010",
    "1111011101001001",
    "1110111110001010",
    "1110100111010101",
    "1110011011001110",
    "1110011010111000",
    "1110100110001110",
    "1110111100001111",
    "1111011010101000",
    "1111111110001110",
    "1111011101010100",
    "1110111101111000",
    "1110101000110100",
    "1110100001010010",
    "1110100111001101",
    "1110110110101010",
    "1111001001100111",
    "1111011001110101",
    "1111100010111001",
    "1111100010111001",
    "1111011100000100",
    "1111010101010000",
    "1111010110001101",
    "1111100010111000",
    "1111111010010110",
    "1111101001000010",
    "1111001110110001",
    "1110111101011001",
    "1110111000111010",
    "1111000000011010",
    "1111001110100011",
    "1111011101101000",
    "1111101011100110",
    "1111111010101110",
    "1111110001111110",
    "1111011010000111",
    "1111000000100001",
    "1110101010110010",
    "1110011111010010",
    "1110100010101100",
    "1110110100110100",
    "1111010000000101",
    "1111101100011001",
    "1111111101111101",
    "1111110011011011",
    "1111110011000000",
    "1111111001010011",
    "1111111111000110",
    "1111111101100000",
    "1111111001100000",
    "1111100101011111",
    "1111001001101010",
    "1110101101001010",
    "1110010110110100",
    "1110001011100011",
    "1110001101101011",
    "1110011010110000",
    "1110101101111111",
    "1111000010010000",
    "1111010010111011",
    "1111100000000000",
    "1111101110001101",
    "1111111110100110",
    "1111100101001000",
    "1111001000010001",
    "1110101111000000",
    "1110011111110011",
    "1110011111010010",
    "1110101110001100",
    "1111000111000001",
    "1111100001010101",
    "1111110101101111",
    "1111111111111001",
    "1111111110110110",
    "1111111100011111",
    "1111110110011001",
    "1111110011010101",
    "1111110110001110",
    "1111111111100001",
    "1111110001111010",
    "1111100001010010",
    "1111010010100010",
    "1111001000001001",
    "1111000011000000",
    "1111000010111101",
    "1111000110111110",
    "1111001101010010",
    "1111010011010111",
    "1111010110011000",
    "1111010100111011",
    "1111001111000101",
    "1111000110000100",
    "1110111011111111",
    "1110110010110001",
    "1110101100100000",
    "1110101100001001",
    "1110110100011100",
    "1111000110001000",
    "1111011111101000",
    "1111111100111010",
    "1111100111010011",
    "1111010010011100",
    "1111001000011011",
    "1111001001101111",
    "1111010011001000",
    "1111100000000000",
    "1111101011101100",
    "1111110010100110",
    "1111110011011100",
    "1111110000011010",
    "1111101110110100",
    "1111110011111011",
    "1111111101111001",
    "1111101000010011",
    "1111010000010010",
    "1110111011111101",
    "1110110000100111",
    "1110110000010100",
    "1110111000101101",
    "1111000101001011",
    "1111010000110001",
    "1111010111011111",
    "1111011000001000",
    "1111010011110001",
    "1111001100111000",
    "1111000110010011",
    "1111000001110001",
    "1110111111010100",
    "1110111110011011",
    "1110111111100110",
    "1111000100100000",
    "1111001110101000",
    "1111011101101110",
    "1111101110111011",
    "1111111101111001",
    "1111111000111010",
    "1111110111000000",
    "1111111010010001",
    "1111111101111010",
    "1111111101001111",
    "1111110101101011",
    "1111100111111001",
    "1111010110111011",
    "1111000110001110",
    "1110111000111010",
    "1110110000110110",
    "1110101110000101",
    "1110101111011010",
    "1110110011011100",
    "1110111000111010",
    "1110111111010111",
    "1111000110011101",
    "1111001101111111",
    "1111010111111110",
    "1111100111010010",
    "1111111101011001",
    "1111100110010000",
    "1111000111100011",
    "1110101100010111",
    "1110011010001100",
    "1110010101001110",
    "1110011101001010",
    "1110101110001001",
    "1111000101110001",
    "1111100010010101",
    "1111111101111110",
    "1111011101000000",
    "1110111110101011",
    "1110100111000001",
    "1110011000101111",
    "1110010101110100",
    "1110011100101011",
    "1110101001000111",
    "1110111001101111",
    "1111001110100110",
    "1111100111101100",
    "1111111011101001",
    "1111011111011111",
    "1111001001010101",
    "1110111110001111",
    "1111000010110110",
    "1111010111010001",
    "1111110110010000",
    "1111100111110000",
    "1111001010111101",
    "1110111001000111",
    "1110110011001101",
    "1110110110010110",
    "1110111101011100",
    "1111000011100001",
    "1111000110010010",
    "1111000110000100",
    "1111000100011100",
    "1111000011110110",
    "1111000111101111",
    "1111010011001011",
    "1111100111001111",
    "1111111101010011",
    "1111011110011100",
    "1111000001011010",
    "1110101011001100",
    "1110011111100110",
    "1110011111011010",
    "1110101000010110",
    "1110110110100101",
    "1111000110011010",
    "1111010100110011",
    "1111100000001000",
    "1111101010000101",
    "1111110110101011",
    "1111110110111010",
    "1111011110101011",
    "1111000100101001",
    "1110101110111111",
    "1110100011011010",
    "1110100101110001",
    "1110110101001011",
    "1111001011110111",
    "1111100100000101",
    "1111111010110011",
    "1111110000001110",
    "1111011011101010",
    "1111000110101100",
    "1110110001111000",
    "1110011110111011",
    "1110010001100001",
    "1110001101111010",
    "1110010111000100",
    "1110101101100100",
    "1111001110111000",
    "1111110101101010",
    "1111100100110001",
    "1111000110011010",
    "1110110010111110",
    "1110101011101011",
    "1110101111001101",
    "1110111010000001",
    "1111000111100010",
    "1111010011011111",
    "1111011011000010",
    "1111011101001110",
    "1111011011000110",
    "1111011001001011",
    "1111011101101000",
    "1111101100000101",
    "1111111011110100",
    "1111011110101101",
    "1111000011011010",
    "1110101111111101",
    "1110101000000011",
    "1110101011011110",
    "1110110110000100",
    "1111000010010111",
    "1111001011100110",
    "1111001111010110",
    "1111001110011011",
    "1111001011001010",
    "1111000111110010",
    "1111000101101110",
    "1111000111000011",
    "1111001110011100",
    "1111011101010100",
    "1111110011000000",
    "1111110011100111",
    "1111011011100000",
    "1111001001010110",
    "1111000001001000",
    "1111000100001110",
    "1111001111101001",
    "1111011101110111",
    "1111101001001010",
    "1111101101110111",
    "1111101011111001",
    "1111100101001011",
    "1111011100011001",
    "1111010100001011",
    "1111001101110101",
    "1111001001001011",
    "1111000101001101",
    "1111000000110011",
    "1110111011100101",
    "1110110110100000",
    "1110110010111101",
    "1110110010000000",
    "1110110011111001",
    "1110111000010000",
    "1111000000011010",
    "1111001111101001",
    "1111100111100010",
    "1111111001001100",
    "1111010110111100",
    "1110111000010011",
    "1110100011001011",
    "1110011011001010",
    "1110011111111010",
    "1110101100000100",
    "1110111000011000",
    "1110111111110011",
    "1111000011100111",
    "1111001001100111",
    "1111010111010001",
    "1111101110101101",
    "1111110010101101",
    "1111010011101111",
    "1110111101100110",
    "1110111010001001",
    "1111001101101001",
    "1111110100001010",
    "1111011100000111",
    "1110101111101000",
    "1110010000001000",
    "1110000001110001",
    "1110000100011101",
    "1110010011001011",
    "1110100110111110",
    "1110111011111111",
    "1111010001101001",
    "1111101000110111",
    "1111111101111000",
    "1111100101011111",
    "1111010010011101",
    "1111001000110100",
    "1111001011000111",
    "1111011000011000",
    "1111101100011101",
    "1111111101010001",
    "1111101001000011",
    "1111011001100010",
    "1111001111000101",
    "1111001001011110",
    "1111001000111001",
    "1111001101110111",
    "1111011001100000",
    "1111101100010011",
    "1111111011100111",
    "1111100001111110",
    "1111001010111000",
    "1110111001100101",
    "1110101110110101",
    "1110101000111110",
    "1110100101001101",
    "1110100000101100",
    "1110011010101011",
    "1110010100100000",
    "1110010001010010",
    "1110010110110110",
    "1110101001111010",
    "1111001011000111",
    "1111110111001001",
    "1111011001101101",
    "1110110000100001",
    "1110010100000011",
    "1110000111111110",
    "1110001010011101",
    "1110010101100100",
    "1110100011010000",
    "1110101110111010",
    "1110110110111111",
    "1110111111001000",
    "1111001100010111",
    "1111100001110100",
    "1111111111010110",
    "1111011111110110",
    "1111000010111001",
    "1110101111110001",
    "1110101010011000",
    "1110110010001101",
    "1111000011000110",
    "1111011000101000",
    "1111101111101100",
    "1111111001100001",
    "1111100011111100",
    "1111010001000111",
    "1111000010110011",
    "1110111010010001",
    "1110111000011101",
    "1110111100111010",
    "1111000101101110",
    "1111010000110101",
    "1111011100101011",
    "1111101001101111",
    "1111111010000110",
    "1111110000100110",
    "1111010110101010",
    "1110111011010100",
    "1110100100001110",
    "1110010111010011",
    "1110011001000100",
    "1110101011010110",
    "1111001011010011",
    "1111110010100000",
    "1111100110011111",
    "1111000110001001",
    "1110110000000000",
    "1110100100111110",
    "1110100100001000",
    "1110101010100110",
    "1110110101100101",
    "1111000011110100",
    "1111010100110011",
    "1111101000001110",
    "1111111100111110",
    "1111101111100010",
    "1111100000000010",
    "1111010101110100",
    "1111010000010111",
    "1111001101010010",
    "1111001001101101",
    "1111000011100010",
    "1110111010000111",
    "1110101110100001",
    "1110100011010011",
    "1110011011010011",
    "1110011000011101",
    "1110011011000001",
    "1110100001100110",
    "1110101010001001",
    "1110110010111000",
    "1110111010011011",
    "1111000000011110",
    "1111000111100011",
    "1111010100000000",
    "1111101000000000",
    "1111111101010001",
    "1111100000000010",
    "1111000110000001",
    "1110110100000000",
    "1110101100101000",
    "1110101111001111",
    "1110110111001000",
    "1110111110111101",
    "1111000101101110",
    "1111001110101011",
    "1111011110001010",
    "1111110101111110",
    "1111101100100110",
    "1111001111010100",
    "1110111000101111",
    "1110101110010001",
    "1110110000100100",
    "1110111011000111",
    "1111001001001011",
    "1111011000100010",
    "1111101000101100",
    "1111111010110000",
    "1111110001011001",
    "1111011111000010",
    "1111010011000110",
    "1111010011100110",
    "1111100011011101",
    "1111111111001001",
    "1111100000111101",
    "1111000110000011",
    "1110110111101101",
    "1110111000100000",
    "1111000101100100",
    "1111011000000110",
    "1111100111111011",
    "1111101111010101",
    "1111101100110100",
    "1111100010010010",
    "1111010100010111",
    "1111001000010101",
    "1111000001110110",
    "1111000010001101",
    "1111001000100101",
    "1111010010100111",
    "1111011101110101",
    "1111100111111001",
    "1111101111000111",
    "1111110100101010",
    "1111111100010001",
    "1111110111011101",
    "1111100110011000",
    "1111010011010010",
    "1111000011001000",
    "1110111010000110",
    "1110111010111100",
    "1111000101100100",
    "1111010101101001",
    "1111100101110001",
    "1111110001000101",
    "1111110101010011",
    "1111110110010010",
    "1111111010011011",
    "1111111001100011",
    "1111100100000110",
    "1111001001001011",
    "1110110000010010",
    "1110100000011001",
    "1110011110100011",
    "1110101010101011",
    "1110111111001101",
    "1111010101001000",
    "1111100110110100",
    "1111110010011011",
    "1111111001100001",
    "1111111111101010",
    "1111110011001111",
    "1111011101001010",
    "1110111110000101",
    "1110011011001001",
    "1101111011111010",
    "1101100111000110",
    "1101100000101011",
    "1101101000010101",
    "1101111001010001",
    "1110001101010111",
    "1110011111100100",
    "1110101100100110",
    "1110110100001110",
    "1110111000000011",
    "1110111010001011",
    "1110111110011100",
    "1111001001111111",
    "1111011111101000",
    "1111111110100010",
    "1111011110000101",
    "1110111110001010",
    "1110101000101100",
    "1110100001101011",
    "1110101001010000",
    "1110111010101011",
    "1111001110101001",
    "1111011110001111",
    "1111100100111110",
    "1111100010100010",
    "1111011010010001",
    "1111010000010100",
    "1111001000100010",
    "1111000100011111",
    "1111000011001111",
    "1111000101011011",
    "1111001110000010",
    "1111011111101000",
    "1111111011001010",
    "1111100001110001",
    "1110111101011110",
    "1110011111011010",
    "1110001110011100",
    "1110001101011001",
    "1110011001000001",
    "1110101010111101",
    "1110111100010100",
    "1111000111101010",
    "1111001101011011",
    "1111010011000000",
    "1111011101111101",
    "1111110001101110",
    "1111110011010001",
    "1111010111100111",
    "1111000010100010",
    "1110111010000100",
    "1110111111101110",
    "1111001110100001",
    "1111011110101011",
    "1111101011011010",
    "1111110100111010",
    "1111111110101111",
    "1111110011110000",
    "1111100010100001",
    "1111010000001101",
    "1111000001001100",
    "1110111010011011",
    "1110111101110011",
    "1111001001100011",
    "1111011100001001",
    "1111110100001011",
    "1111110000011011",
    "1111010011101111",
    "1110111001100011",
    "1110100110110100",
    "1110011111101011",
    "1110100111101100",
    "1110111111110000",
    "1111100100011100",
    "1111110000011100",
    "1111000110111111",
    "1110100110101100",
    "1110010100000101",
    "1110010000100111",
    "1110011010001110",
    "1110101011111101",
    "1111000000101011",
    "1111010011100111",
    "1111100001001100",
    "1111100111111011",
    "1111101000010101",
    "1111100100011000",
    "1111011111000100",
    "1111011011011011",
    "1111011011110010",
    "1111100000111000",
    "1111101001100111",
    "1111110011100011",
    "1111111100010000",
    "1111111101001010",
    "1111110111011110",
    "1111110000100001",
    "1111100111001110",
    "1111011100001110",
    "1111010001011010",
    "1111001001011011",
    "1111000110010101",
    "1111001000100011",
    "1111001110100011",
    "1111010100111011",
    "1111010111111111",
    "1111010101101001",
    "1111001110011001",
    "1111000101001000",
    "1110111101011100",
    "1110111010001100",
    "1110111100010110",
    "1111000011001010",
    "1111001100100001",
    "1111010101101010",
    "1111011101000010",
    "1111100100001011",
    "1111101101110101",
    "1111111011011000",
    "1111110011101111",
    "1111100010010010",
    "1111010011101001",
    "1111001010110100",
    "1111001001100011",
    "1111001110111000",
    "1111010111011011",
    "1111011111011010",
    "1111100011110110",
    "1111100011011010",
    "1111011110011100",
    "1111010111100010",
    "1111010100100010",
    "1111011011000001",
    "1111101100110100",
    "1111111000011110",
    "1111011011011000",
    "1111000011011100",
    "1110110110011010",
    "1110110110110010",
    "1111000010000000",
    "1111010010010000",
    "1111100001010101",
    "1111101010111010",
    "1111110000010010",
    "1111110110101000",
    "1111111101100111",
    "1111101010011010",
    "1111010001110011",
    "1110111001011101",
    "1110100111001101",
    "1110011111011001",
    "1110100010010010",
    "1110101011110010",
    "1110110110100101",
    "1110111110010100",
    "1111000011111110",
    "1111001101100001",
    "1111011111111111",
    "1111111100111101",
    "1111011110010110",
    "1110111001001100",
    "1110011011011001",
    "1110001011000111",
    "1110001010100010",
    "1110010101111100",
    "1110100110011011",
    "1110110101011010",
    "1110111111001000",
    "1111000011111011",
    "1111000110100000",
    "1111001001111010",
    "1111010000011110",
    "1111011001110111",
    "1111100011000011",
    "1111101000010110",
    "1111100110101000",
    "1111011100110111",
    "1111001101010001",
    "1110111100100001",
    "1110101111010111",
    "1110101001001100",
    "1110101011100000",
    "1110110101101111",
    "1111000101110010",
    "1111010111111001",
    "1111101000100101",
    "1111111000010110",
    "1111110101111000",
    "1111100000000011",
    "1111000110000000",
    "1110101010100101",
    "1110010010011010",
    "1110000010000101",
    "1101111101100001",
    "1110000101001000",
    "1110010101001001",
    "1110101000100000",
    "1110111010001011",
    "1111000111010101",
    "1111001111100011",
    "1111010011011111",
    "1111010111010101",
    "1111100001001111",
    "1111110100011010",
    "1111101111101010",
    "1111001111111011",
    "1110110011111110",
    "1110100010011100",
    "1110011111001111",
    "1110101001101011",
    "1110111100011100",
    "1111010001010100",
    "1111100010100110",
    "1111101100100000",
    "1111101111000110",
    "1111101100110101",
    "1111101001001100",
    "1111101000101100",
    "1111101111111100",
    "1111111110101111",
    "1111100100010010",
    "1111000100111100",
    "1110100111011011",
    "1110010001011110",
    "1110000110010110",
    "1110000110110111",
    "1110010000001101",
    "1110011101100000",
    "1110101010010001",
    "1110110100101010",
    "1110111110111101",
    "1111001101010100",
    "1111100010001011",
    "1111111100111010",
    "1111100110101111",
    "1111001110110110",
    "1110111111110110",
    "1110111010111101",
    "1110111101101011",
    "1111000011000001",
    "1111000110001101",
    "1111000100110111",
    "1111000000000111",
    "1110111010111111",
    "1110111000100000",
    "1110111010000100",
    "1110111111101011",
    "1111001001010000",
    "1111010111001011",
    "1111101001110110",
    "1111111111001101",
    "1111100101100100",
    "1111001011010100",
    "1110110011010011",
    "1110100000110101",
    "1110010110011000",
    "1110010100000101",
    "1110010111101010",
    "1110011101101001",
    "1110100010110011",
    "1110100100110001",
    "1110100100101100",
    "1110100111011011",
    "1110110001110110",
    "1111000110100000",
    "1111100011011000",
    "1111111101100111",
    "1111100011011100",
    "1111010011100001",
    "1111001111101100",
    "1111010100100010",
    "1111011100100110",
    "1111100010101110",
    "1111100011101110",
    "1111011111111111",
    "1111011001101111",
    "1111010100010111",
    "1111010100000011",
    "1111011010101011",
    "1111100110110111",
    "1111110100100011",
    "1111111101100100",
    "1111111100010000",
    "1111101110011110",
    "1111010110011000",
    "1110111010001110",
    "1110100001101110",
    "1110010011001010",
    "1110010001110001",
    "1110011100100101",
    "1110101110101101",
    "1111000011000101",
    "1111011000001000",
    "1111101110111001",
    "1111110110011101",
    "1111010111000011",
    "1110110101010011",
    "1110010101110010",
    "1101111101111010",
    "1101110010000000",
    "1101110010010101",
    "1101111011010011",
    "1110000111111010",
    "1110010011111000",
    "1110011101011100",
    "1110100101100101",
    "1110101101100100",
    "1110110111110111",
    "1111001000101101",
    "1111100010111110",
    "1111111001110000",
    "1111010001011100",
    "1110101010111101",
    "1110001101010001",
    "1101111101010110",
    "1101111101011100",
    "1110001011001110",
    "1110100000110110",
    "1110111000000110",
    "1111001011000111",
    "1111010111101101",
    "1111100001100111",
    "1111101110011110",
    "1111111101100011",
    "1111100001111000",
    "1111000011001000",
    "1110101000000011",
    "1110010110101100",
    "1110010010111101",
    "1110011011110111",
    "1110101110010001",
    "1111000111010001",
    "1111100011101010",
    "1111111111000011",
    "1111100011110100",
    "1111001110001111",
    "1111000000101001",
    "1110111011110011",
    "1110111111111000",
    "1111001100111000",
    "1111100010111110",
    "1111111111000110",
    "1111011101000100",
    "1110111100010110",
    "1110100010111001",
    "1110010100110110",
    "1110010100101001",
    "1110100011001101",
    "1110111110101001",
    "1111100010010010",
    "1111111000010101",
    "1111010111100000",
    "1110111111100100",
    "1110110010111000",
    "1110110000010100",
    "1110110100000110",
    "1110111010110111",
    "1111000010101001",
    "1111001011011101",
    "1111010110001001",
    "1111100010110001",
    "1111101111011100",
    "1111111001111001",
    "1111111111010001",
    "1111111100010011",
    "1111111100000101",
    "1111111100101001",
    "1111111011011111",
    "1111110110010101",
    "1111101100010101",
    "1111011110111010",
    "1111010001100100",
    "1111001000010000",
    "1111000101100010",
    "1111001001100000",
    "1111010010010111",
    "1111011101010001",
    "1111100110111011",
    "1111101100101011",
    "1111101101000101",
    "1111101000001100",
    "1111011111110000",
    "1111010110111100",
    "1111010011000011",
    "1111011001011101",
    "1111101100010101",
    "1111110110011110",
    "1111010100101001",
    "1110110101000011",
    "1110011101011001",
    "1110010001001100",
    "1110010000110000",
    "1110011001000001",
    "1110100101101110",
    "1110110011010000",
    "1110111111110011",
    "1111001011111010",
    "1111011001001001",
    "1111101000101001",
    "1111111010001011",
    "1111110100111001",
    "1111101000010011",
    "1111100010111110",
    "1111100110001000",
    "1111110000100111",
    "1111111111010010",
    "1111110001101101",
    "1111100100111100",
    "1111011010111101",
    "1111010011000110",
    "1111001100010100",
    "1111000101101110",
    "1110111110101110",
    "1110110111101101",
    "1110110001110001",
    "1110101110010100",
    "1110110000010001",
    "1110111011001111",
    "1111010001000011",
    "1111110000100010",
    "1111101010101101",
    "1111000111101000",
    "1110101101000101",
    "1110100000010001",
    "1110100010100100",
    "1110110000101011",
    "1111000100011111",
    "1111010111100010",
    "1111100110111100",
    "1111110101001110",
    "1111111001111000",
    "1111100100011101",
    "1111001011110011",
    "1110110101010000",
    "1110100111000110",
    "1110100110000001",
    "1110110010110100",
    "1111001000100101",
    "1111011111010001",
    "1111101111011101",
    "1111110100111110",
    "1111110000011100",
    "1111100101101111",
    "1111011001011110",
    "1111010001100010",
    "1111010011010000",
    "1111100000010010",
    "1111110110110001",
    "1111101110010011",
    "1111010101110001",
    "1111000100101111",
    "1110111101111000",
    "1111000001001000",
    "1111001011001010",
    "1111010111010001",
    "1111100001000111",
    "1111100101101010",
    "1111100100110100",
    "1111100000010001",
    "1111011001101101",
    "1111010011001101",
    "1111001110001100",
    "1111001010100011",
    "1111001000001110",
    "1111001001100000",
    "1111010001111101",
    "1111100011111011",
    "1111111110110011",
    "1111100010001000",
    "1111000110010011",
    "1110110100100111",
    "1110110001100010",
    "1110111100101101",
    "1111010010001010",
    "1111101110010100",
    "1111110010001111",
    "1111010011001111",
    "1110110111100000",
    "1110100010100001",
    "1110010110111011",
    "1110010110011010",
    "1110100010000011",
    "1110110111110010",
    "1111010010001000",
    "1111101010101010",
    "1111111011010101",
    "1111111111000111",
    "1111111011101101",
    "1111101111100000",
    "1111100010001010",
    "1111011001011101",
    "1111011001001001",
    "1111100011001011",
    "1111110110101110",
    "1111101111110001",
    "1111010100111011",
    "1110111101100100",
    "1110101110010010",
    "1110101010011011",
    "1110110010011111",
    "1111000011011100",
    "1111010111111100",
    "1111101010011111",
    "1111110111011000",
    "1111111110011100",
    "1111111101110000",
    "1111111010001011",
    "1111110100011010",
    "1111101100000100",
    "1111100010110011",
    "1111011011101000",
    "1111011001011001",
    "1111011100110111",
    "1111100011111011",
    "1111101011001001",
    "1111101111100010",
    "1111101111101110",
    "1111101100011110",
    "1111101001100010",
    "1111101100110100",
    "1111111010100000",
    "1111101101011010",
    "1111001111100001",
    "1110110011010111",
    "1110100000011110",
    "1110011100000010",
    "1110100110101100",
    "1110111011011110",
    "1111010010110110",
    "1111100101101010",
    "1111101110111111",
    "1111101101100110",
    "1111100011011000",
    "1111010011101111",
    "1111000010110001",
    "1110110011101110",
    "1110101000011010",
    "1110100001101110",
    "1110011111100011",
    "1110100001111101",
    "1110101010100000",
    "1110111010111000",
    "1111010010111011",
    "1111101111100111",
    "1111110011110100",
    "1111011011110000",
    "1111001011000110",
    "1111000010110100",
    "1111000001010101",
    "1111000011011000",
    "1111000101011011",
    "1111000100110001",
    "1111000000100111",
    "1110111001110100",
    "1110110010000101",
    "1110101011011110",
    "1110101000000110",
    "1110101011001111",
    "1110111000001001",
    "1111001111101100",
    "1111101111101100",
    "1111101100110111",
    "1111001100011011",
    "1110110100101111",
    "1110101001111010",
    "1110101101001111",
    "1110111101110111",
    "1111011001001011",
    "1111111011011100",
    "1111011111111000",
    "1110111101111000",
    "1110100011111011",
    "1110010110011101",
    "1110010111011011",
    "1110100101001110",
    "1110111010101010",
    "1111010001110001",
    "1111100111100001",
    "1111111011110110",
    "1111110000010001",
    "1111011100010111",
    "1111001001010000",
    "1110111001001110",
    "1110101111011100",
    "1110101110101101",
    "1110110110110110",
    "1111000100001000",
    "1111010001100111",
    "1111011010110000",
    "1111011110111010",
    "1111100011010011",
    "1111101101110001",
    "1111111110011110",
    "1111100010011111",
    "1111000100010010",
    "1110101011101000",
    "1110011111000010",
    "1110100001100111",
    "1110110000011100",
    "1111000101000101",
    "1111011001000111",
    "1111101000001001",
    "1111110011011101",
    "1111111111110011",
    "1111101111101101",
    "1111011010100101",
    "1111000100000001",
    "1110110010010111",
    "1110101010110010",
    "1110101111111010",
    "1110111111110110",
    "1111010011110100",
    "1111100100100000",
    "1111101101001000",
    "1111101100110001",
    "1111100110001011",
    "1111011101000100",
    "1111010100110011",
    "1111010001111110",
    "1111011000101101",
    "1111101010000101",
    "1111111011011011",
    "1111011100100101",
    "1111000000000010",
    "1110101011011110",
    "1110100010111101",
    "1110100111011000",
    "1110110101100010",
    "1111001010010100",
    "1111100011011000",
    "1111111110001101",
    "1111100110110011",
    "1111001110100011",
    "1110111100101101",
    "1110110011011000",
    "1110110100000110",
    "1110111110010010",
    "1111001110000101",
    "1111011111010100",
    "1111110000001001",
    "1111111110101011",
    "1111101011001111",
    "1111010100100111",
    "1110111100001100",
    "1110100101010011",
    "1110010100101010",
    "1110001110010010",
    "1110010010011100",
    "1110011101101011",
    "1110101010111101",
    "1110110101111001",
    "1110111100011110",
    "1111000000001000",
    "1111000110001011",
    "1111010100111110",
    "1111101111011110",
    "1111101100100010",
    "1111000110001000",
    "1110100110001101",
    "1110010100000101",
    "1110010011010101",
    "1110100010010000",
    "1110111010001001",
    "1111010011100100",
    "1111101001000011",
    "1111110111110110",
    "1111111111110110",
    "1111111110100110",
    "1111111100110011",
    "1111110010111100",
    "1111100100011111",
    "1111010011000000",
    "1111000001110011",
    "1110110101101110",
    "1110110100010101",
    "1111000001000010",
    "1111011010101000",
    "1111111011110001",
    "1111100010111011",
    "1111000111101101",
    "1110110101101010",
    "1110101100101101",
    "1110101010011000",
    "1110101011011101",
    "1110101101101001",
    "1110101111110000",
    "1110110001011001",
    "1110110010101001",
    "1110110011111011",
    "1110110110100100",
    "1110111101000010",
    "1111001001100010",
    "1111011100100001",
    "1111110100000100",
    "1111110011001111",
    "1111011101000111",
    "1111001100100001",
    "1111000011101010",
    "1111000100000001",
    "1111001110000101",
    "1111100000111001",
    "1111111010100011",
    "1111100111101011",
    "1111001001100011",
    "1110101111011111",
    "1110011110000100",
    "1110011000100111",
    "1110100001110000",
    "1110111010110101",
    "1111100010000101",
    "1111101101111011",
    "1110111101010001",
    "1110010100110110",
    "1101111011110111",
    "1101110110000011",
    "1110000010101001",
    "1110011100000010",
    "1110111010010011",
    "1111010101110100",
    "1111101001100001",
    "1111110011110000",
    "1111110111001010",
    "1111111010110111",
    "1111111001101111",
    "1111100011101010",
    "1111000101001101",
    "1110100101010111",
    "1110001100100000",
    "1110000001010111",
    "1110000111010101",
    "1110011011101000",
    "1110111000001000",
    "1111011001000110",
    "1111111101001010",
    "1111011100010001",
    "1110110100001101",
    "1110001110011111",
    "1101110000001101",
    "1101011110001001",
    "1101011100111100",
    "1101101100101110",
    "1110001000100000",
    "1110101001001110",
    "1111000110110111",
    "1111011100001111",
    "1111101011000111",
    "1111111000111011",
    "1111110100100011",
    "1111011010110000",
    "1110111100110111",
    "1110100001001111",
    "1110001101110011",
    "1110000110111011",
    "1110001011110111",
    "1110010111000100",
    "1110100010100100",
    "1110101010000110",
    "1110101100110010",
    "1110101100111000",
    "1110101100110010",
    "1110101110010001",
    "1110110100101100",
    "1111000011001111",
    "1111011010011000",
    "1111111000000110",
    "1111101000011010",
    "1111001100110010",
    "1110111001011000",
    "1110110001010000",
    "1110110100101110",
    "1110111111111111",
    "1111001101010110",
    "1111010110111001",
    "1111011000101111",
    "1111010010110100",
    "1111000111101100",
    "1110111011001111",
    "1110110001110000",
    "1110101100111111",
    "1110101100100001",
    "1110101110110101",
    "1110110001101110",
    "1110110011101010",
    "1110110100110011",
    "1110111000010000",
    "1111000010100001",
    "1111010110000110",
    "1111110010100011",
    "1111101011100011",
    "1111001010010110",
    "1110110000001101",
    "1110100001100110",
    "1110011110110110",
    "1110100011101111",
    "1110101010100110",
    "1110101110111000",
    "1110101110010111",
    "1110101010000001",
    "1110100100011010",
    "1110100010010100",
    "1110101001111111",
    "1110111110100011",
    "1111011110111010",
    "1111111010000001",
    "1111010100000001",
    "1110110110000000",
    "1110100100100000",
    "1110100000101100",
    "1110100111001001",
    "1110110011010111",
    "1111000010111011",
    "1111010101011000",
    "1111101011011110",
    "1111111010110011",
    "1111100000000011",
    "1111001000011000",
    "1110111000101010",
    "1110110101100100",
    "1111000000100100",
    "1111010111011010",
    "1111110101000011",
    "1111101101011010",
    "1111010110100100",
    "1111001010000001",
    "1111001000010000",
    "1111001111000010",
    "1111011010100110",
    "1111100110111001",
    "1111110000001011",
    "1111110100001010",
    "1111110011000111",
    "1111101111000010",
    "1111101010101010",
    "1111101000011111",
    "1111101010101010",
    "1111110011010011",
    "1111111100111011",
    "1111101000001000",
    "1111010010001101",
    "1111000000000111",
    "1110110110010101",
    "1110110111110111",
    "1111000101100010",
    "1111011101010111",
    "1111111011001110",
    "1111100101001110",
    "1111000111111010",
    "1110101111101110",
    "1110011110010110",
    "1110010100101111",
    "1110010011011101",
    "1110011010010110",
    "1110101000011010",
    "1110111011010001",
    "1111001111101001",
    "1111100010010010",
    "1111110001011111",
    "1111111111000011",
    "1111110000111110",
    "1111011011010100",
    "1110111111010110",
    "1110100000110001",
    "1110000110110001",
    "1101111010100011",
    "1110000011110011",
    "1110100011100111",
    "1111010011111000",
    "1111110110001001",
    "1111000111000100",
    "1110101010000110",
    "1110100101100101",
    "1110111000111111",
    "1111011100011011",
    "1111111011101001",
    "1111011001110100",
    "1111000100100100",
    "1110111101001111",
    "1111000000010111",
    "1111000111110100",
    "1111001110000101",
    "1111010010100010",
    "1111011001100111",
    "1111101000001101",
    "1111111111001001",
    "1111011110100001",
    "1110111100011001",
    "1110100000111101",
    "1110010010111011",
    "1110010100111110",
    "1110100011101001",
    "1110111000001001",
    "1111001011100110",
    "1111011001010001",
    "1111100001101100",
    "1111101010001101",
    "1111111000011110",
    "1111101111111011",
    "1111001111111101",
    "1110101101000010",
    "1110001101111101",
    "1101111001000010",
    "1101110010001010",
    "1101111000011011",
    "1110000111010011",
    "1110011001100010",
    "1110101010101101",
    "1110111000110100",
    "1111000011010101",
    "1111001011101101",
    "1111010110100101",
    "1111101000011000",
    "1111111101110000",
    "1111011110001100",
    "1110111110011111",
    "1110100101001000",
    "1110010110111110",
    "1110010110001001",
    "1110100000010100",
    "1110110000000010",
    "1110111111101001",
    "1111001010011011",
    "1111001110011100",
    "1111001100110101",
    "1111001000011011",
    "1111000100110110",
    "1111000100111100",
    "1111001001101010",
    "1111010010111101",
    "1111011111110001",
    "1111101110100011",
    "1111111110000101",
    "1111110010010000",
    "1111100010100111",
    "1111010011011000",
    "1111000101010111",
    "1110111001000111",
    "1110101110110110",
    "1110100110101100",
    "1110100001000101",
    "1110011110100100",
    "1110011111000010",
    "1110100001101100",
    "1110100101100010",
    "1110101010000100",
    "1110101111001000",
    "1110110100110011",
    "1110111011000110",
    "1111000001110000",
    "1111001000011101",
    "1111001110011001",
    "1111010011011000",
    "1111011001100000",
    "1111100100011101",
    "1111110110101000",
    "1111110000000101",
    "1111010010111101",
    "1110110111000100",
    "1110100001011001",
    "1110010101100101",
    "1110010100100101",
    "1110011100000101",
    "1110101000010000",
    "1110110101000110",
    "1110111111101100",
    "1111000111110100",
    "1111001111010001",
    "1111011000110111",
    "1111100111011000",
    "1111111100000010",
    "1111101001110011",
    "1111001100110011",
    "1110110001011010",
    "1110011100000111",
    "1110001111111011",
    "1110001101101001",
    "1110010100001011",
    "1110100001010100",
    "1110110001110000",
    "1111000010010100",
    "1111010011001000",
    "1111100110110111",
    "1111111111110000",
    "1111100001111110",
    "1111000001110001",
    "1110100101011000",
    "1110010010010000",
    "1110001011111010",
    "1110010001111000",
    "1110011111000010",
    "1110101100110101",
    "1110110111110101",
    "1111000001011100",
    "1111001101001111",
    "1111011101111101",
    "1111110011011101",
    "1111110101010100",
    "1111100001011010",
    "1111010101110111",
    "1111010101000110",
    "1111011100111101",
    "1111101010100011",
    "1111111100100110",
    "1111101101111111",
    "1111010101110001",
    "1110111100100110",
    "1110100110101010",
    "1110011000010000",
    "1110010101110010",
    "1110100001001111",
    "1110110111010000",
    "1111010001111110",
    "1111101011010110",
    "1111111110010011",
    "1111110111010100",
    "1111110101011100",
    "1111111010001111",
    "1111111101011000",
    "1111110100010110",
    "1111101100111011",
    "1111101001011101",
    "1111101010111001",
    "1111110000010010",
    "1111110111101001",
    "1111111110011010",
    "1111111110001111",
    "1111111110100001",
    "1111110010101110",
    "1111011110101000",
    "1111000100101111",
    "1110101001010001",
    "1110010001011001",
    "1110000001101110",
    "1101111101001111",
    "1110000100001101",
    "1110010011111001",
    "1110100111101101",
    "1110111011000010",
    "1111001010010110",
    "1111010100010011",
    "1111011001100000",
    "1111011011011110",
    "1111011011101101",
    "1111011100110010",
    "1111100010110110",
    "1111110001010011",
    "1111110110111110",
    "1111011000011110",
    "1110111000100101",
    "1110011101010110",
    "1110001100000111",
    "1110000111111001",
    "1110001111000010",
    "1110011100100000",
    "1110101010100101",
    "1110110101000001",
    "1110111010011101",
    "1110111011101011",
    "1110111100010100",
    "1111000010011100",
    "1111010010011001",
    "1111101100001111",
    "1111110011101100",
    "1111010100000101",
    "1110111011001001",
    "1110101101010111",
    "1110101011111101",
    "1110110011110110",
    "1111000000010100",
    "1111001100111010",
    "1111010110010110",
    "1111011100000100",
    "1111011111000111",
    "1111100001001111",
    "1111100100011111",
    "1111101001011010",
    "1111101110111011",
    "1111110011100001",
    "1111110101100100",
    "1111110100000100",
    "1111101111010010",
    "1111101000100011",
    "1111100001101001",
    "1111011011111000",
    "1111011000011011",
    "1111011000001000",
    "1111011100000001",
    "1111100110000011",
    "1111110111101100",
    "1111101111100011",
    "1111010010010000",
    "1110110100101100",
    "1110011011111100",
    "1110001100010110",
    "1110001000011110",
    "1110001111011111",
    "1110011101001110",
    "1110101100010110",
    "1110111000010000",
    "1110111110001100",
    "1110111110100001",
    "1110111101000101",
    "1110111111100001",
    "1111001010011101",
    "1111011110111000",
    "1111111001010011",
    "1111101100100101",
    "1111011001100011",
    "1111010010001010",
    "1111010110011111",
    "1111100001111101",
    "1111101110011100",
    "1111110110111011",
    "1111111001000110",
    "1111110110000001",
    "1111110000101001",
    "1111101100010001",
    "1111101011001110",
    "1111101101101001",
    "1111110010000001",
    "1111110110001001",
    "1111111000001011",
    "1111110111100000",
    "1111110100100100",
    "1111110010100101",
    "1111110110111001",
    "1111111011000100",
    "1111100011010011",
    "1111000101011011",
    "1110101000000110",
    "1110010001111001",
    "1110000111110010",
    "1110001011100001",
    "1110011001100011",
    "1110101011110101",
    "1110111100011011",
    "1111000111011111",
    "1111001111011001",
    "1111011001111101",
    "1111101011100001",
    "1111111010010010",
    "1111011011010011",
    "1110111111000111",
    "1110101100111100",
    "1110101010000010",
    "1110110110110110",
    "1111001101101011",
    "1111100110110101",
    "1111111011100011",
    "1111110110111001",
    "1111101101011000",
    "1111100010101001",
    "1111010010011010",
    "1110111010110000",
    "1110011110010111",
    "1110000011010011",
    "1101101111111111",
    "1101101001011000",
    "1101110000001101",
    "1110000000101001",
    "1110010101000101",
    "1110101000101101",
    "1110111010111010",
    "1111001110001111",
    "1111100100101010",
    "1111111110011110",
    "1111100110011000",
    "1111001110011111",
    "1110111110011111",
    "1110111001011110",
    "1110111111101110",
    "1111001110100001",
    "1111100010011100",
    "1111111000001100",
    "1111110011010000",
    "1111100010110001",
    "1111011001101000",
    "1111011011001010",
    "1111101001000101",
    "1111111101100100",
    "1111011101001010",
    "1110111100101010",
    "1110100010111001",
    "1110010100001110",
    "1110010001011010",
    "1110010111100111",
    "1110100001111101",
    "1110101100001010",
    "1110110100001010",
    "1110111010010011",
    "1111000000010101",
    "1111000111011010",
    "1111010000100011",
    "1111011110010110",
    "1111110011001000",
    "1111110000101001",
    "1111001110101110",
    "1110101011011000",
    "1110001100000111",
    "1101110110010000",
    "1101101110001101",
    "1101110100011100",
    "1110000101001011",
    "1110011011000111",
    "1110110000011111",
    "1111000001010000",
    "1111001011110011",
    "1111010010001111",
    "1111011010100011",
    "1111101010011011",
    "1111111100000111",
    "1111011011110010",
    "1110111011001100",
    "1110100001111001",
    "1110010101101111",
    "1110011000100000",
    "1110100111100101",
    "1110111111000101",
    "1111011011010100",
    "1111111000100110",
    "1111101011100001",
    "1111010010111110",
    "1110111111000111",
    "1110110000111000",
    "1110101001000111",
    "1110101000001100",
    "1110101110000000",
    "1110111010110101",
    "1111001110100100",
    "1111100111110011",
    "1111111100010011",
    "1111100001010111",
    "1111001010101111",
    "1110111011011001",
    "1110110110010101",
    "1110111101101000",
    "1111010001001000",
    "1111101101111111",
    "1111110000110101",
    "1111010001010010",
    "1110111000010110",
    "1110101000111110",
    "1110100100000110",
    "1110101000110100",
    "1110110100101100",
    "1111000110101100",
    "1111011111000010",
    "1111111101011111",
    "1111011111100001",
    "1110111011110111",
    "1110011100101010",
    "1110000110100010",
    "1101111100110000",
    "1101111111011110",
    "1110001010110101",
    "1110011001101111",
    "1110100111001001",
    "1110110000110110",
    "1110111010011101",
    "1111001010000100",
    "1111100011101110",
    "1111111000110000",
    "1111010001011110",
    "1110101111000000",
    "1110011000101000",
    "1110010011000001",
    "1110011101000010",
    "1110110000010001",
    "1111000100110110",
    "1111010101000011",
    "1111100001100110",
    "1111110000000111",
    "1111111011001010",
    "1111011111010010",
    "1110111111110110",
    "1110100100011111",
    "1110010100100010",
    "1110010100101001",
    "1110100100001000",
    "1110111100001001",
    "1111010011111100",
    "1111100100011111",
    "1111101010110100",
    "1111101000110010",
    "1111100001101001",
    "1111011000010101",
    "1111001111000100",
    "1111000110001101",
    "1110111101000000",
    "1110110011001111",
    "1110101010100101",
    "1110100111100011",
    "1110101110110110",
    "1111000001111011",
    "1111011101010110",
    "1111111001110010",
    "1111110000010111",
    "1111100110001011",
    "1111101000011100",
    "1111110011101000",
    "1111111110001011",
    "1111110010100100",
    "1111101100100000",
    "1111101011110001",
    "1111101110011010",
    "1111110010011000",
    "1111110110000101",
    "1111111000010100",
    "1111111000000010",
    "1111110100011110",
    "1111101101001000",
    "1111100010011100",
    "1111010101101001",
    "1111001001011000",
    "1111000010100100",
    "1111000111001001",
    "1111011010001100",
    "1111111010000011",
    "1111011111111111",
    "1110111101010100",
    "1110100101111011",
    "1110011110011110",
    "1110100110111100",
    "1110111010001111",
    "1111010001010010",
    "1111100101011000",
    "1111110010010010",
    "1111110111001000",
    "1111110101010001",
    "1111101110101111",
    "1111100110101111",
    "1111100000111000",
    "1111011111110011",
    "1111100100011100",
    "1111101101110000",
    "1111111001110011",
    "1111111001010011",
    "1111101101110011",
    "1111100101110110",
    "1111100010011010",
    "1111100010111001",
    "1111100101011010",
    "1111100111110001",
    "1111101000011011",
    "1111100110101101",
    "1111100010100010",
    "1111011101100100",
    "1111011100001001",
    "1111100010110011",
    "1111110011011111",
    "1111110011010101",
    "1111010111001001",
    "1110111110010010",
    "1110101101101011",
    "1110100111111001",
    "1110101011100101",
    "1110110011111100",
    "1110111011110000",
    "1110111111010001",
    "1110111101111111",
    "1110111100101110",
    "1111000010011111",
    "1111010100010011",
    "1111110011000101",
    "1111100110010000",
    "1111000000110000",
    "1110100101010010",
    "1110011010101010",
    "1110100010010010",
    "1110110110111100",
    "1111010000010111",
    "1111100111000011",
    "1111111000000101",
    "1111111001110111",
    "1111101011001011",
    "1111011001101101",
    "1111000101100111",
    "1110110010101111",
    "1110100110011011",
    "1110100100111001",
    "1110101111011110",
    "1111000010111011",
    "1111011001111100",
    "1111110000111001",
    "1111111001000011",
    "1111100010111000",
    "1111001011011110",
    "1110110011110110",
    "1110011110110101",
    "1110010000100110",
    "1110001111001101",
    "1110011111110011",
    "1111000010110100",
    "1111110011110100",
    "1111010110000100",
    "1110100101100000",
    "1110000010110100",
    "1101110010011111",
    "1101110100000110",
    "1110000010010100",
    "1110010101111100",
    "1110101000111010",
    "1110111001110101",
    "1111001101000000",
    "1111100110101010",
    "1111111000000111",
    "1111010010001010",
    "1110101101111000",
    "1110010001111101",
    "1110000011101001",
    "1110000100100111",
    "1110010001001010",
    "1110100010110001",
    "1110110011100111",
    "1111000010001010",
    "1111010010000101",
    "1111100111010111",
    "1111111100111100",
    "1111011100111010",
    "1110111101110011",
    "1110100101101010",
    "1110011001000110",
    "1110011001111010",
    "1110100101110110",
    "1110110111100101",
    "1111001001100010",
    "1111010111110111",
    "1111100001011110",
    "1111100110111111",
    "1111101011001011",
    "1111110010011101",
    "1111111111101100",
    "1111101100111111",
    "1111010110011111",
    "1111000001100110",
    "1110110011000000",
    "1110101110000000",
    "1110110011001011",
    "1110111111110000",
    "1111010000010111",
    "1111100010111001",
    "1111110110000010",
    "1111110110111101",
    "1111100101100000",
    "1111010111111111",
    "1111010000101001",
    "1111010000110101",
    "1111011000010011",
    "1111100100100000",
    "1111110001011110",
    "1111111100000010",
    "1111111101010111",
    "1111111010111100",
    "1111111011011100",
    "1111111101011111",
    "1111111110110010",
    "1111111011111110",
    "1111110011000001",
    "1111100011110100",
    "1111001111111101",
    "1110111011001001",
    "1110101001110101",
    "1110100000000111",
    "1110100000011100",
    "1110101001101010",
    "1110111000010000",
    "1111000111111100",
    "1111010100101001",
    "1111011100000010",
    "1111011110000000",
    "1111011101001111",
    "1111011111000010",
    "1111100111100100",
    "1111110111101000",
    "1111110011011111",
    "1111011111001101",
    "1111010001010010",
    "1111001101100100",
    "1111010100100010",
    "1111100010111001",
    "1111110011100101",
    "1111111101110011",
    "1111110011011010",
    "1111101100010001",
    "1111100101010101",
    "1111011011010100",
    "1111001100100110",
    "1110111010010100",
    "1110101000011101",
    "1110011011111010",
    "1110011000000011",
    "1110011101010001",
    "1110101000111010",
    "1110110110100010",
    "1111000001110100",
    "1111001000011000",
    "1111001010100000",
    "1111001100000001",
    "1111010010101011",
    "1111100010110100",
    "1111111101100000",
    "1111100000100011",
    "1110111110000000",
    "1110100010000011",
    "1110010010010010",
    "1110010000001111",
    "1110011000110000",
    "1110100110010110",
    "1110110011100100",
    "1110111100111010",
    "1111000001111110",
    "1111000100001011",
    "1111000101100000",
    "1111001000000001",
    "1111001110010111",
    "1111011011011000",
    "1111110000000101",
    "1111110101001111",
    "1111011001000001",
    "1111000000101100",
    "1110110000110110",
    "1110101100101101",
    "1110110100010010",
    "1111000011011100",
    "1111010100100000",
    "1111100010010101",
    "1111101010000011",
    "1111101011101001",
    "1111101001010000",
    "1111101000001011",
    "1111101110100000",
    "1111111110110100",
    "1111101000010111",
    "1111001101010110",
    "1110111001110100",
    "1110110110100000",
    "1111000111110001",
    "1111101011001000",
    "1111101000111000",
    "1110111111111000",
    "1110100100000001",
    "1110011100110111",
    "1110101100101000",
    "1111001111111010",
    "1111111111000111",
    "1111001111110000",
    "1110100101101010",
    "1110001000001011",
    "1101111001110010",
    "1101111001000111",
    "1110000001010010",
    "1110001101011001",
    "1110011010110000",
    "1110101001000001",
    "1110111001001100",
    "1111001011010100",
    "1111011101011001",
    "1111101100001110",
    "1111110100010001",
    "1111110011010010",
    "1111101010010000",
    "1111011101001110",
    "1111010001111101",
    "1111001111010001",
    "1111011010001011",
    "1111110010110110",
    "1111101011010101",
    "1111001000011110",
    "1110101100111010",
    "1110011110010001",
    "1110011110101110",
    "1110101100100101",
    "1111000010001010",
    "1111011000100000",
    "1111101010001000",
    "1111110100000000",
    "1111110110000111",
    "1111110010111100",
    "1111101111011001",
    "1111110001010001",
    "1111111011110000",
    "1111110010000111",
    "1111011100100110",
    "1111001001011001",
    "1110111101011100",
    "1110111011000110",
    "1111000001101011",
    "1111001110001010",
    "1111011101100000",
    "1111101101111010",
    "1111111110111000",
    "1111101111101010",
    "1111011110010111",
    "1111001110111111",
    "1111000100000110",
    "1111000000110000",
    "1111000111001110",
    "1111010111110100",
    "1111110000110001",
    "1111110001011111",
    "1111010011101110",
    "1110111010110101",
    "1110101010011110",
    "1110100011110100",
    "1110100101110110",
    "1110101101111101",
    "1110111000110111",
    "1111000011000101",
    "1111001010110100",
    "1111010010001111",
    "1111011101011100",
    "1111101111011011",
    "1111110111110000",
    "1111011011110010",
    "1111000010001000",
    "1110110000001000",
    "1110101001011000",
    "1110101101011110",
    "1110111000101100",
    "1111000111011010",
    "1111011000001000",
    "1111101011110011",
    "1111111011110011",
    "1111011111011001",
    "1111000010001011",
    "1110101001010101",
    "1110011010101010",
    "1110011010010011",
    "1110101000111001",
    "1111000100000110",
    "1111100111100111",
    "1111110001101000",
    "1111001011111111",
    "1110101010110000",
    "1110010000100111",
    "1101111111110101",
    "1101111001111010",
    "1101111110110110",
    "1110001100010100",
    "1110011110011100",
    "1110110001111000",
    "1111000110001011",
    "1111011101000111",
    "1111111000000010",
    "1111101001010101",
    "1111001010000100",
    "1110101111000111",
    "1110011101101001",
    "1110011001001011",
    "1110100000110000",
    "1110101111000101",
    "1110111101101001",
    "1111000111000011",
    "1111001000110101",
    "1111000110011011",
    "1111000111001000",
    "1111010001100001",
    "1111101000001011",
    "1111111000101000",
    "1111011001100101",
    "1111000101110100",
    "1111000111101101",
    "1111100010100010",
    "1111110000001011",
    "1110111101011110",
    "1110010011011101",
    "1101111100011011",
    "1101111100001001",
    "1110001111100011",
    "1110101110010111",
    "1111010001010000",
    "1111110101000100",
    "1111100111000011",
    "1111000011001011",
    "1110100001001100",
    "1110000101000000",
    "1101110010110110",
    "1101101110011111",
    "1101111000001110",
    "1110001011010001",
    "1110100001010111",
    "1110110101001011",
    "1111000011101111",
    "1111001100111111",
    "1111010010010111",
    "1111010101111110",
    "1111011011010001",
    "1111100110001110",
    "1111111001000011",
    "1111101100100011",
    "1111001110000111",
    "1110110001010111",
    "1110011011110111",
    "1110010010001010",
    "1110010110011111",
    "1110100110100101",
    "1110111100111111",
    "1111010011001000",
    "1111100011001010",
    "1111101001111111",
    "1111100111101011",
    "1111011110011100",
    "1111010010110011",
    "1111001010010011",
    "1111001001001001",
    "1111010000111101",
    "1111011111100001",
    "1111101111100011",
    "1111111011100101",
    "1111111111111001",
    "1111111100011101",
    "1111110011111100",
    "1111101100101001",
    "1111101100101010",
    "1111110110111100",
    "1111110110100111",
    "1111100001111001",
    "1111010001010100",
    "1111001001110010",
    "1111001101001111",
    "1111011001110111",
    "1111101011101110",
    "1111111110100010",
    "1111110001000100",
    "1111100100110111",
    "1111011101000010",
    "1111011000100000",
    "1111010101110100",
    "1111010011111011",
    "1111010010000000",
    "1111001111010100",
    "1111001011111010",
    "1111001000100111",
    "1111000110101100",
    "1111000111011011",
    "1111001011101101",
    "1111010100110100",
    "1111100100100100",
    "1111111011101110",
    "1111100110111110",
    "1111000110101101",
    "1110100111110010",
    "1110001110011111",
    "1101111101110111",
    "1101110110110100",
    "1101110111111110",
    "1101111110000010",
    "1110000101011000",
    "1110001011100110",
    "1110010000001010",
    "1110010011101110",
    "1110010111111111",
    "1110100000000101",
    "1110101111010001",
    "1111000110100101",
    "1111100100000110",
    "1111111101000011",
    "1111100011011010",
    "1111010100110110",
    "1111010101000000",
    "1111100011011101",
    "1111111011100110",
    "1111101001011101",
    "1111010010100001",
    "1111000100001010",
    "1110111111001111",
    "1111000010000000",
    "1111001010010100",
    "1111010111100111",
    "1111101010010011",
    "1111111101100001",
    "1111100001010100",
    "1111000100000110",
    "1110101010001100",
    "1110011000010000",
    "1110010001011100",
    "1110010101111001",
    "1110100010110011",
    "1110110100010111",
    "1111001001001001",
    "1111100010101100",
    "1111111101100001",
    "1111011000000110",
    "1110110000100011",
    "1110001101000100",
    "1101110100000011",
    "1101101010010011",
    "1101110000101110",
    "1110000010111101",
    "1110011001110100",
    "1110101110100001",
    "1110111100110101",
    "1111000100101111",
    "1111001000110010",
    "1111001011111000",
    "1111010010101001",
    "1111100010000011",
    "1111111100000000",
    "1111100001001100",
    "1110111011000100",
    "1110011001010000",
    "1110000001111011",
    "1101111001000110",
    "1101111111101011",
    "1110010001110100",
    "1110101001000010",
    "1110111110100011",
    "1111001100110010",
    "1111010010110110",
    "1111010101011000",
    "1111011010101111",
    "1111101000001010",
    "1111111110111101",
    "1111100100111011",
    "1111001001111111",
    "1110110110101000",
    "1110101111010100",
    "1110110011001000",
    "1110111100111000",
    "1111000110110111",
    "1111001101000010",
    "1111001110010010",
    "1111001100001001",
    "1111001000101100",
    "1111000110101010",
    "1111001000111010",
    "1111010000111000",
    "1111011110101001",
    "1111110000100111",
    "1111111100000011",
    "1111101010010111",
    "1111011100101010",
    "1111010100111110",
    "1111010100011111",
    "1111011010110111",
    "1111100101101100",
    "1111110001001110",
    "1111111001100110",
    "1111111011110010",
    "1111110110001010",
    "1111101000110010",
    "1111010101010111",
    "1110111110100001",
    "1110100111100111",
    "1110010100000110",
    "1110000111000110",
    "1110000011000001",
    "1110001001110101",
    "1110011100000100",
    "1110110111111110",
    "1111011001010011",
    "1111111010100100",
    "1111101001000100",
    "1111010100101111",
    "1111001001000100",
    "1111000011111110",
    "1111000001110001",
    "1110111110111111",
    "1110111010001100",
    "1110110100011100",
    "1110110000000111",
    "1110101111011100",
    "1110110011100100",
    "1110111100010110",
    "1111001000111111",
    "1111011001011011",
    "1111101110001100",
    "1111111000101000",
    "1111011100010011",
    "1110111111010100",
    "1110100101100111",
    "1110010100000000",
    "1110001110011111",
    "1110010110101111",
    "1110101011000010",
    "1111000111010000",
    "1111100110000011",
    "1111111101111010",
    "1111101001001100",
    "1111011110101011",
    "1111011111101011",
    "1111101100000110",
    "1111111101010110",
    "1111011111011110",
    "1110111110110011",
    "1110100001001000",
    "1110001100000001",
    "1110000011010000",
    "1110000111100000",
    "1110010110001110",
    "1110101010100010",
    "1110111110111101",
    "1111001111010010",
    "1111011001100010",
    "1111011110010010",
    "1111100001001100",
    "1111100111001101",
    "1111110100000100",
    "1111110111101100",
    "1111011111010100",
    "1111001000001000",
    "1110110111100010",
    "1110110001101110",
    "1110111000010011",
    "1111001001110010",
    "1111100010111001",
    "1111111111111100",
    "1111100010011001",
    "1111000111001110",
    "1110110001110110",
    "1110100101100100",
    "1110100100100111",
    "1110101111110001",
    "1111000101110100",
    "1111100011001011",
    "1111111101011110",
    "1111100010000101",
    "1111001111001010",
    "1111000110001101",
    "1111000101000011",
    "1111000111001110",
    "1111001000010001",
    "1111000101101100",
    "1110111111100011",
    "1110110111101111",
    "1110110000110110",
    "1110101100111000",
    "1110101110010001",
    "1110111000011110",
    "1111001101100000",
    "1111101100011000",
    "1111101110110001",
    "1111001010100101",
    "1110101101100100",
    "1110011100110000",
    "1110011011101011",
    "1110101011111101",
    "1111001011111000",
    "1111110110101001",
    "1111011011001110",
    "1110110010001111",
    "1110010101011000",
    "1110001001000001",
    "1110001101010110",
    "1110011101111011",
    "1110110100011000",
    "1111001100110000",
    "1111100111001000",
    "1111111011000010",
    "1111011001101011",
    "1110111000000001",
    "1110011011001111",
    "1110001000010000",
    "1110000011001101",
    "1110001101000000",
    "1110100001011100",
    "1110111001101000",
    "1111001110101101",
    "1111011100001010",
    "1111100010001000",
    "1111100011111011",
    "1111100111000111",
    "1111110001111111",
    "1111111000100011",
    "1111011010100101",
    "1110111001011011",
    "1110011100100000",
    "1110001010000110",
    "1110000101110010",
    "1110001111110001",
    "1110100100011101",
    "1110111110001111",
    "1111010111011010",
    "1111101011010101",
    "1111110111101000",
    "1111111100001111",
    "1111111010101001",
    "1111110101000001",
    "1111101101100010",
    "1111100101100111",
    "1111011110111101",
    "1111011100011110",
    "1111100001001000",
    "1111101110011101",
    "1111111100011011",
    "1111100010111110",
    "1111001010000010",
    "1110110110011111",
    "1110101011100101",
    "1110101001111010",
    "1110101111011100",
    "1110111000110000",
    "1111000010011001",
    "1111001001110101",
    "1111001110101001",
    "1111010010100110",
    "1111011000101101",
    "1111100011100110",
    "1111110011100100",
    "1111111001111000",
    "1111101001000011",
    "1111011110001101",
    "1111011011110010",
    "1111100000110110",
    "1111101010000000",
    "1111110011010101",
    "1111111001111100",
    "1111111101000000",
    "1111111101110011",
    "1111111110100011",
    "1111111110110000",
    "1111111001101011",
    "1111110011100100",
    "1111101110101111",
    "1111101101000000",
    "1111101110111110",
    "1111110011100111",
    "1111111000110000",
    "1111111100001101",
    "1111111100101011",
    "1111111001101010",
    "1111110011000011",
    "1111101000110101",
    "1111011011100000",
    "1111001100100101",
    "1110111110110101",
    "1110110110001101",
    "1110110110101000",
    "1111000010101110",
    "1111011010001001",
    "1111111001011101",
    "1111100100110001",
    "1111000110000100",
    "1110101110100110",
    "1110100000001101",
    "1110011010010110",
    "1110011010110000",
    "1110011110101000",
    "1110100011101010",
    "1110101000110101",
    "1110101101110000",
    "1110110010001000",
    "1110110101101010",
    "1110111000000001",
    "1110111001000010",
    "1110111001000010",
    "1110111000101111",
    "1110111001001100",
    "1110111100000010",
    "1111000011000110",
    "1111001111010110",
    "1111011111111000",
    "1111110001110100",
    "1111111111010110",
    "1111111000010000",
    "1111111011100001",
    "1111110111010100",
    "1111100100010111",
    "1111010001110000",
    "1111000101010010",
    "1111000011111000",
    "1111010001010010",
    "1111101101101011",
    "1111101011000011",
    "1111000000001101",
    "1110011010011110",
    "1110000001000010",
    "1101110111111001",
    "1101111111010100",
    "1110010010101011",
    "1110101010110111",
    "1111000001011111",
    "1111010010000011",
    "1111011101011001",
    "1111101001000100",
    "1111111010000100",
    "1111101100111101",
    "1111001110000010",
    "1110101111110001",
    "1110011001010110",
    "1110010000011111",
    "1110010111010000",
    "1110101001100011",
    "1111000000000111",
    "1111010100001011",
    "1111100001100111",
    "1111101000001000",
    "1111101001011111",
    "1111100111111100",
    "1111100101101110",
    "1111100101001000",
    "1111101001011011",
    "1111110101011001",
    "1111110110111001",
    "1111011110011011",
    "1111000110001011",
    "1110110011011111",
    "1110101010011101",
    "1110101100101011",
    "1110110111010110",
    "1111000100010101",
    "1111001101011011",
    "1111001110110011",
    "1111001000011110",
    "1110111101100001",
    "1110110010010000",
    "1110101010110000",
    "1110101010011001",
    "1110110011011010",
    "1111000110000001",
    "1111100000000111",
    "1111111101010011",
    "1111100111101000",
    "1111010011001011",
    "1111001000010000",
    "1111000111101101",
    "1111001110111010",
    "1111011001000100",
    "1111100001100001",
    "1111100101011111",
    "1111100100111011",
    "1111100001010111",
    "1111011100100110",
    "1111011000001100",
    "1111010100101100",
    "1111010001101110",
    "1111001110111010",
    "1111001100001111",
    "1111001010100000",
    "1111001010111111",
    "1111001110110101",
    "1111010110000100",
    "1111100000100111",
    "1111101111100110",
    "1111111011101101",
    "1111100001110011",
    "1111000101011010",
    "1110101011001110",
    "1110011000000011",
    "1110001111000111",
    "1110010001011001",
    "1110011100001111",
    "1110101010011011",
    "1110110110110100",
    "1110111101111011",
    "1110111111101001",
    "1111000000001111",
    "1111000101011111",
    "1111010011001011",
    "1111101000110100",
    "1111111110101011",
    "1111101010011011",
    "1111100000011001",
    "1111100011101110",
    "1111110010110011",
    "1111111000000101",
    "1111100011011100",
    "1111010100000011",
    "1111001100001010",
    "1111001011100110",
    "1111010001010010",
    "1111011011011011",
    "1111100111111101",
    "1111110101010010",
    "1111111101100100",
    "1111110001010011",
    "1111100101111001",
    "1111011011011110",
    "1111010010100111",
    "1111001100001010",
    "1111001001011101",
    "1111001100000101",
    "1111010101011011",
    "1111100110000110",
    "1111111100111101",
    "1111101001000001",
    "1111010000010100",
    "1110111101100011",
    "1110110011111001",
    "1110110011111001",
    "1110111011111111",
    "1111001010000010",
    "1111011100110010",
    "1111110011100011",
    "1111110010011011",
    "1111010110100100",
    "1110111011000100",
    "1110100011001000",
    "1110010010001010",
    "1110001010100010",
    "1110001100100101",
    "1110010110101100",
    "1110100101110100",
    "1110110110011000",
    "1111000101011010",
    "1111010001001010",
    "1111011011001100",
    "1111101000100011",
    "1111111101100110",
    "1111100100101111",
    "1111000001111011",
    "1110100000111001",
    "1110001000110101",
    "1101111110101110",
    "1110000100010011",
    "1110010101111100",
    "1110101101000101",
    "1111000110001110",
    "1111100001000010",
    "1111111110100010",
    "1111100001000010",
    "1111000000111001",
    "1110100110010101",
    "1110010110011111",
    "1110010101101001",
    "1110100011010111",
    "1110111001110010",
    "1111010001000111",
    "1111100001110001",
    "1111100111100001",
    "1111100010110011",
    "1111011000001100",
    "1111001111111000",
    "1111010001101100",
    "1111100000011001",
    "1111111001100111",
    "1111101001000011",
    "1111001111101110",
    "1111000000100111",
    "1110111110100001",
    "1111000111010101",
    "1111010101100010",
    "1111100011011000",
    "1111101101111111",
    "1111110111100000",
    "1111111011101011",
    "1111101000110110",
    "1111010000000111",
    "1110110101100101",
    "1110011111011110",
    "1110010011100010",
    "1110010100110110",
    "1110100001011110",
    "1110110011100111",
    "1111000100110100",
    "1111010000000000",
    "1111010011011111",
    "1111010000010101",
    "1111001010000001",
    "1111000111000001",
    "1111001101100110",
    "1111100000011111",
    "1111111110000111",
    "1111011111100011",
    "1111000000100110",
    "1110101100000010",
    "1110100110001000",
    "1110101110001010",
    "1110111111010111",
    "1111010011100100",
    "1111100100110001",
    "1111101111010101",
    "1111110010100011",
    "1111101111101011",
    "1111101001010101",
    "1111100010011111",
    "1111011100010001",
    "1111010101110001",
    "1111001101000010",
    "1111000000100111",
    "1110110001100111",
    "1110100100101111",
    "1110100000100111",
    "1110101010000010",
    "1111000001100111",
    "1111100011010101",
    "1111111000011100",
    "1111011010011000",
    "1111001001001110",
    "1111000110111110",
    "1111010000000000",
    "1111011101001010",
    "1111100110111011",
    "1111101000100010",
    "1111100001100010",
    "1111010110010000",
    "1111001110110110",
    "1111010010101110",
    "1111100100011101",
    "1111111110101100",
    "1111011110000010",
    "1111000001111000",
    "1110110000111011",
    "1110101110000000",
    "1110110110101101",
    "1111000101010011",
    "1111010011111110",
    "1111011111111011",
    "1111101011100000",
    "1111111010111010",
    "1111101111000111",
    "1111010011000101",
    "1110110101110110",
    "1110011110110101",
    "1110010100100100",
    "1110011010000111",
    "1110101100101000",
    "1111000100111001",
    "1111011010100010",
    "1111100111101001",
    "1111101101010000",
    "1111110000111101",
    "1111111000010010",
    "1111111001100101",
    "1111100110001000",
    "1111010010100010",
    "1111000100111100",
    "1111000010000110",
    "1111001010110010",
    "1111011010110101",
    "1111101100110010",
    "1111111110010111",
    "1111101111010001",
    "1111011010011110",
    "1111000011010010",
    "1110101100101101",
    "1110011011000111",
    "1110010011000000",
    "1110010111100010",
    "1110100111100111",
    "1110111111110001",
    "1111011110010010",
    "1111111110100000",
    "1111011000101000",
    "1110110010010000",
    "1110010000001101",
    "1101110111111111",
    "1101101101111111",
    "1101110101000001",
    "1110001010010100",
    "1110101000011101",
    "1111001100001010",
    "1111110010010100",
    "1111100111100010",
    "1111000011011100",
    "1110100100001101",
    "1110001100000100",
    "1101111101100110",
    "1101111100001001",
    "1110001000011110",
    "1110100001101110",
    "1111000101010000",
    "1111101101110111",
    "1111101001111110",
    "1111000111011111",
    "1110101110010111",
    "1110011111011110",
    "1110011001011000",
    "1110011001101101",
    "1110011101100110",
    "1110100011011111",
    "1110101100000010",
    "1110111001000010",
    "1111001100000001",
    "1111100101001000",
    "1111111101011100",
    "1111011111110001",
    "1111000110100101",
    "1110110101101010",
    "1110101110010001",
    "1110101110111011",
    "1110110100110110",
    "1110111100110111",
    "1111000101001001",
    "1111001101100011",
    "1111010110011101",
    "1111100000001111",
    "1111101010100110",
    "1111110011111100",
    "1111111001101010",
    "1111111001000101",
    "1111110000100100",
    "1111100000010001",
    "1111001010010100",
    "1110110010101001",
    "1110011101111010",
    "1110001111101100",
    "1110001001100101",
    "1110001011001100",
    "1110010011011000",
    "1110100000111011",
    "1110110010100111",
    "1111000111110100",
    "1111011111111010",
    "1111111010000001",
    "1111101010111010",
    "1111010000011010",
    "1110111000001001",
    "1110100011110011",
    "1110010100110001",
    "1110001011110011",
    "1110001000101000",
    "1110001010001111",
    "1110001111010001",
    "1110010101110110",
    "1110011100011100",
    "1110100010000011",
    "1110100110001110",
    "1110101001010001",
    "1110101011101010",
    "1110101111101000",
    "1110111001010011",
    "1111001011000100",
    "1111100100001110",
    "1111111110110011",
    "1111100011111000",
    "1111010000000011",
    "1111000110101010",
    "1111000111111111",
    "1111010000001100",
    "1111011001101000",
    "1111011111100011",
    "1111011111001000",
    "1111011000110111",
    "1111001111010110",
    "1111000101011010",
    "1110111101111000",
    "1110111010001110",
    "1110111010000100",
    "1110111100100001",
    "1111000000011111",
    "1111000101010010",
    "1111001010110100",
    "1111010001000111",
    "1111010111110010",
    "1111011101110010",
    "1111100010000011",
    "1111100100010000",
    "1111100101001000",
    "1111100101100010",
    "1111100110110100",
    "1111101100001011",
    "1111111001100011",
    "1111101111000100",
    "1111001110111111",
    "1110101011010001",
    "1110001010111111",
    "1101110100011101",
    "1101101100001001",
    "1101110010100001",
    "1110000011100110",
    "1110011001010011",
    "1110101101111000",
    "1110111101011110",
    "1111000111011010",
    "1111001100010011",
    "1111001110110011",
    "1111010100101100",
    "1111100010101011",
    "1111111001110000",
    "1111101000110000",
    "1111001011011011",
    "1110110110101101",
    "1110110010110110",
    "1111000100100101",
    "1111101001111000",
    "1111100101100101",
    "1110110100111100",
    "1110001110101101",
    "1101111001010011",
    "1101110101001110",
    "1101111101111011",
    "1110001100010001",
    "1110011011101101",
    "1110101101010110",
    "1111000100010101",
    "1111100010100001",
    "1111111001100000",
    "1111010101010101",
    "1110111000011101",
    "1110101010001100",
    "1110101111010010",
    "1111000111011011",
    "1111101101110111",
    "1111100101010000",
    "1110111011100011",
    "1110011100111101",
    "1110001101110000",
    "1110001111001100",
    "1110011111000000",
    "1110111000101000",
    "1111010110111100",
    "1111110100111010",
    "1111110001100011",
    "1111011111000101",
    "1111010101000011",
    "1111010011010111",
    "1111010111111110",
    "1111011111100011",
    "1111100110110000",
    "1111101011001000",
    "1111101100000010",
    "1111101010001100",
    "1111100111000011",
    "1111100100011100",
    "1111100011111000",
    "1111100110010011",
    "1111101011101111",
    "1111110011001000",
    "1111111011001011",
    "1111111100111001",
    "1111110101100110",
    "1111101110111011",
    "1111101001000011",
    "1111100100100101",
    "1111100001111001",
    "1111100000011111",
    "1111011110111111",
    "1111011011011001",
    "1111010100110001",
    "1111001011100000",
    "1111000001011100",
    "1110111001010001",
    "1110110101001011",
    "1110110110110111",
    "1111000001001010",
    "1111010110010010",
    "1111110101111000",
    "1111100011001011",
    "1110111011100001",
    "1110011010011110",
    "1110000101100010",
    "1101111111101000",
    "1110000111001101",
    "1110010110111001",
    "1110101000010011",
    "1110110101110100",
    "1110111100100101",
    "1110111101000000",
    "1110111000111111",
    "1110110011010000",
    "1110101110010010",
    "1110101011001010",
    "1110101010010011",
    "1110101100100110",
    "1110110011111110",
    "1111000010100111",
    "1111011001011000",
    "1111110110100010",
    "1111101010000111",
    "1111001110010010",
    "1110111011000001",
    "1110110010100001",
    "1110110011101110",
    "1110111011000001",
    "1111000011111011",
    "1111001010100101",
    "1111001100110101",
    "1111001010001001",
    "1111000011100110",
    "1110111011011000",
    "1110110011101001",
    "1110101101111101",
    "1110101011001111",
    "1110101100000100",
    "1110110000110101",
    "1110111001110101",
    "1111001000000001",
    "1111011101001001",
    "1111111001101100",
    "1111100100010111",
    "1111000001001111",
    "1110100010010010",
    "1110001100101010",
    "1110000011110100",
    "1110001000101101",
    "1110011000100010",
    "1110101101101000",
    "1111000001110110",
    "1111010000010100",
    "1111010110101101",
    "1111010101011000",
    "1111001110100110",
    "1111000101110100",
    "1110111110011001",
    "1110111010100011",
    "1110111011001110",
    "1110111111101001",
    "1111000101100111",
    "1111001010011011",
    "1111001011111100",
    "1111001001011001",
    "1111000011011100",
    "1110111100000100",
    "1110110110000011",
    "1110110011111110",
    "1110111001000001",
    "1111001000110010",
    "1111100100000101",
    "1111110111110100",
    "1111010000111011",
    "1110101111000010",
    "1110011000101101",
    "1110010001110001",
    "1110011001111001",
    "1110101100001001",
    "1111000001110001",
    "1111010101000000",
    "1111100100101110",
    "1111110100111111",
    "1111110110000010",
    "1111011011011110",
    "1110111110010010",
    "1110100101000011",
    "1110010110010101",
    "1110010110010000",
    "1110100100100101",
    "1110111011100000",
    "1111010010111000",
    "1111100100001101",
    "1111101100101000",
    "1111101110001001",
    "1111101100101100",
    "1111101100100001",
    "1111110010000110",
    "1111111111110110",
    "1111101011000000",
    "1111010001101001",
    "1110111000101111",
    "1110100101000001",
    "1110011010000001",
    "1110011001010110",
    "1110100010010111",
    "1110110010100110",
    "1111000110001110",
    "1111011001000001",
    "1111100111010100",
    "1111101111010001",
    "1111110010101100",
    "1111110110100010",
    "1111111111101000",
    "1111101111110001",
    "1111011001001100",
    "1111000001010111",
    "1110101110010001",
    "1110100100110111",
    "1110100110110001",
    "1110110000111011",
    "1110111110111111",
    "1111001110011111",
    "1111011111001010",
    "1111110001111110",
    "1111111000000000",
    "1111011111010110",
    "1111000101111011",
    "1110101111011010",
    "1110100000011010",
    "1110011100100001",
    "1110100101111011",
    "1110111011111100",
    "1111011010100011",
    "1111111011011101",
    "1111101000001000",
    "1111010101101111",
    "1111010000010100",
    "1111010111100111",
    "1111100111101000",
    "1111111001111100",
    "1111110110010011",
    "1111101001010011",
    "1111011100001001",
    "1111001100000001",
    "1110111000000110",
    "1110100010101110",
    "1110010000011001",
    "1110000110100101",
    "1110001001100000",
    "1110011000011110",
    "1110101110011001",
    "1111000110110110",
    "1111100000101011",
    "1111111101000000",
    "1111100010011101",
    "1110111110101110",
    "1110011011110010",
    "1101111110111111",
    "1101101110011011",
    "1101101101110011",
    "1101111011011110",
    "1110010010001111",
    "1110101011011011",
    "1111000001001100",
    "1111010000110110",
    "1111011010101101",
    "1111100000111011",
    "1111100110001011",
    "1111101100011100",
    "1111110110010101",
    "1111111001011110",
    "1111100010110001",
    "1111000111111001",
    "1110101101011100",
    "1110011000100101",
    "1110001101011011",
    "1110001110011100",
    "1110011010101000",
    "1110101100111111",
    "1110111111001100",
    "1111001100000101",
    "1111010001110000",
    "1111010001010111",
    "1111001101101011",
    "1111001001111010",
    "1111001001101011",
    "1111010000011111",
    "1111100000011111",
    "1111111001001011",
    "1111101000111100",
    "1111001010101000",
    "1110101111110101",
    "1110011011001010",
    "1110001110011011",
    "1110001001101010",
    "1110001011010100",
    "1110010001101001",
    "1110011011001010",
    "1110100111010001",
    "1110110101100010",
    "1111000100101010",
    "1111010011001011",
    "1111011111111010",
    "1111101100011001",
    "1111111100011001",
    "1111101101101111",
    "1111010010010101",
    "1110110100100010",
    "1110011001101011",
    "1110000111000001",
    "1110000000110110",
    "1110000111110010",
    "1110010111011011",
    "1110101001100000",
    "1110111000101101",
    "1111000001111001",
    "1111000101001000",
    "1111000101110110",
    "1111001010011110",
    "1111011000100011",
    "1111110001001000",
    "1111101111111100",
    "1111010010000010",
    "1110111100011110",
    "1110110011111100",
    "1110111000001000",
    "1111000011010101",
    "1111001110010110",
    "1111010011011111",
    "1111010000000111",
    "1111000101101001",
    "1110110111110001",
    "1110101011110010",
    "1110101000111010",
    "1110110100010000",
    "1111001110000101",
    "1111110010100011",
    "1111100110001011",
    "1111000100101110",
    "1110101111011001",
    "1110101001000100",
    "1110101111011110",
    "1110111100101010",
    "1111001010000111",
    "1111010010100001",
    "1111010011010011",
    "1111001101111111",
    "1111001000001000",
    "1111001000100011",
    "1111010011001000",
    "1111100110010010",
    "1111111100010111",
    "1111110001010000",
    "1111100111111101",
    "1111101010000011",
    "1111110101011110",
    "1111111010110101",
    "1111101100001100",
    "1111100010100010",
    "1111100000000101",
    "1111100101010111",
    "1111110001110111",
    "1111111011111111",
    "1111100101110010",
    "1111001100010100",
    "1110110000110110",
    "1110010101110010",
    "1101111110010100",
    "1101101110000010",
    "1101100111110010",
    "1101101100100011",
    "1101111010100101",
    "1110001101111111",
    "1110100010110110",
    "1110111000011011",
    "1111010001000000",
    "1111101110100111",
    "1111101110101101",
    "1111001010010001",
    "1110101010001100",
    "1110010101000110",
    "1110010000001101",
    "1110011101010100",
    "1110111000111001",
    "1111011011110111",
    "1111111110001101",
    "1111100110110000",
    "1111010110001101",
    "1111010000001101",
    "1111010100100100",
    "1111100010100111",
    "1111111001000101",
    "1111101010011011",
    "1111001100010001",
    "1110110001100111",
    "1110011110111111",
    "1110010111011111",
    "1110011011000010",
    "1110100110000001",
    "1110110011011101",
    "1111000000000011",
    "1111001101000000",
    "1111011110010110",
    "1111110110101101",
    "1111101010001000",
    "1111000111111010",
    "1110101000111111",
    "1110010011110001",
    "1110001100100001",
    "1110010010111001",
    "1110100001111110",
    "1110110011011111",
    "1111000010001111",
    "1111001100011110",
    "1111010011100001",
    "1111011010110101",
    "1111101000000100",
    "1111111111001101",
    "1111100000010111",
    "1110111011110011",
    "1110011011000001",
    "1110000101100000",
    "1101111111100001",
    "1110001001000001",
    "1110011101011011",
    "1110110101110111",
    "1111001100010111",
    "1111011100110111",
    "1111100101110010",
    "1111101000110001",
    "1111101010111111",
    "1111110010110111",
    "1111111100000011",
    "1111100011000101",
    "1111000111011011",
    "1110110000011001",
    "1110100100000001",
    "1110100101100100",
    "1110110100111011",
    "1111001111110001",
    "1111110010010011",
    "1111101000001100",
    "1111000100111001",
    "1110101000110000",
    "1110010111100000",
    "1110010100011000",
    "1110100010011010",
    "1111000000111101",
    "1111101011010011",
    "1111100110000011",
    "1110111100101010",
    "1110100000001101",
    "1110010101011101",
    "1110011101010010",
    "1110110010001000",
    "1111001011011001",
    "1111100010010000",
    "1111110010010101",
    "1111111011000001",
    "1111111110100000",
    "1111111111011101",
    "1111111010010010",
    "1111101111000100",
    "1111011101110011",
    "1111001000110000",
    "1110110100000011",
    "1110100100001011",
    "1110011100000100",
    "1110011100010100",
    "1110100011000101",
    "1110101101111010",
    "1110111010110000",
    "1111001000001000",
    "1111010100110011",
    "1111011111011111",
    "1111100111011011",
    "1111101100011010",
    "1111101110010001",
    "1111101101000000",
    "1111101010011101",
    "1111101010111110",
    "1111110010010101",
    "1111111110001100",
    "1111101000010101",
    "1111010000110101",
    "1110111101100000",
    "1110110011001101",
    "1110110100000101",
    "1110111101100011",
    "1111001010011110",
    "1111010110011011",
    "1111011110001101",
    "1111100001010100",
    "1111100010011100",
    "1111100101101010",
    "1111101110101001",
    "1111111110010001",
    "1111101110100100",
    "1111011101001110",
    "1111010010111011",
    "1111010011000011",
    "1111011101001100",
    "1111101101011000",
    "1111111110101000",
    "1111110010101001",
    "1111101000011100",
    "1111100011011010",
    "1111100011010011",
    "1111100111000010",
    "1111101100101010",
    "1111110001111010",
    "1111110100011111",
    "1111110010011111",
    "1111101011001011",
    "1111011111010110",
    "1111010001000101",
    "1111000011101111",
    "1110111010111111",
    "1110111001010011",
    "1110111111000111",
    "1111001001111100",
    "1111010110001000",
    "1111100010010111",
    "1111101111111011",
    "1111111111000010",
    "1111101001011110",
    "1111010001001101",
    "1110111010101011",
    "1110101010110101",
    "1110100101100111",
    "1110101011001111",
    "1110110111100000",
    "1111000100101001",
    "1111001101110000",
    "1111010000011110",
    "1111001110011011",
    "1111001100011001",
    "1111010000010111",
    "1111011110100001",
    "1111110110001000",
    "1111101101111011",
    "1111010100010010",
    "1111000010001011",
    "1110111001111010",
    "1110111001101111",
    "1110111101011100",
    "1111000001001100",
    "1111000011011100",
    "1111000100111001",
    "1111000111000011",
    "1111001010100110",
    "1111001111001111",
    "1111010011101110",
    "1111010110001000",
    "1111010100101100",
    "1111001110110110",
    "1111000101011111",
    "1110111010100101",
    "1110110000011111",
    "1110101001011001",
    "1110100110010011",
    "1110100110100000",
    "1110101000011010",
    "1110101010101010",
    "1110101100011100",
    "1110101101101101",
    "1110101110101101",
    "1110101111111101",
    "1110110010011101",
    "1110110111000110",
    "1111000000001111",
    "1111010001110001",
    "1111101101110000",
    "1111101100111011",
    "1111000011000110",
    "1110011100010110",
    "1101111111110000",
    "1101110010010100",
    "1101110101100101",
    "1110000101101010",
    "1110011011110101",
    "1110110001010111",
    "1111000001011111",
    "1111001100101010",
    "1111010111101111",
    "1111100110111111",
    "1111111100000101",
    "1111101011111001",
    "1111010111111100",
    "1111001110011100",
    "1111010011001111",
    "1111100101011101",
    "1111111110011010",
    "1111101010110011",
    "1111011101010100",
    "1111011100000111",
    "1111100101000110",
    "1111110011101000",
    "1111111101000110",
    "1111110001100001",
    "1111101011101000",
    "1111101010110101",
    "1111101101011010",
    "1111110000111111",
    "1111110011100001",
    "1111110100110100",
    "1111110101111001",
    "1111111000001000",
    "1111111100010111",
    "1111111101011100",
    "1111110110001000",
    "1111101110110010",
    "1111101000110101",
    "1111100101001001",
    "1111100011101001",
    "1111100011100010",
    "1111100011101010",
    "1111100011001101",
    "1111100010000110",
    "1111100001000111",
    "1111100001100110",
    "1111100100111110",
    "1111101011111101",
    "1111110110000110",
    "1111111110001111",
    "1111110011100111",
    "1111101100110100",
    "1111101100101000",
    "1111110100100100",
    "1111111100000111",
    "1111101000111010",
    "1111010110110110",
    "1111001010110000",
    "1111000111100111",
    "1111001101010111",
    "1111011001001100",
    "1111100110100000",
    "1111110000101001",
    "1111110100001011",
    "1111101111101010",
    "1111100011010101",
    "1111010000110101",
    "1110111011001100",
    "1110100110000011",
    "1110010100110100",
    "1110001010000111",
    "1110000111010001",
    "1110001011110101",
    "1110010101110001",
    "1110100010000011",
    "1110101111001101",
    "1110111110101110",
    "1111010010100111",
    "1111101011011110",
    "1111111000010010",
    "1111011101010001",
    "1111001000101000",
    "1110111110010100",
    "1110111111100001",
    "1111001001000010",
    "1111010100111110",
    "1111011101101101",
    "1111011111100110",
    "1111011010100110",
    "1111010001100001",
    "1111000111110100",
    "1111000000110001",
    "1110111110001101",
    "1111000000001000",
    "1111000111011000",
    "1111010101010000",
    "1111101001110011",
    "1111111100010101",
    "1111100000100011",
    "1111000111101000",
    "1110110110100000",
    "1110110000101011",
    "1110110110111111",
    "1111000111101100",
    "1111011111011001",
    "1111111001101100",
    "1111101101111111",
    "1111011011010001",
    "1111010000011010",
    "1111001110001100",
    "1111010011011000",
    "1111011101010110",
    "1111101000100010",
    "1111110010011000",
    "1111111011000101",
    "1111111011000011",
    "1111101110001011",
    "1111011110000000",
    "1111001100001001",
    "1110111011100101",
    "1110110000111000",
    "1110110001111110",
    "1111000010101111",
    "1111100010100010",
    "1111110011101100",
    "1111001000011010",
    "1110100100010011",
    "1110001101110000",
    "1110000111010101",
    "1110001110101011",
    "1110011111100100",
    "1110110111100011",
    "1111010100110001",
    "1111110101101000",
    "1111101000000111",
    "1111001000100101",
    "1110101111101001",
    "1110100000110110",
    "1110100000010101",
    "1110110000001111",
    "1111001110101001",
    "1111110110110111",
    "1111011110110001",
    "1110111010011001",
    "1110100001101100",
    "1110011001100011",
    "1110100100100000",
    "1111000000011001",
    "1111101000001000",
    "1111101100000101",
    "1111000101010111",
    "1110101010000100",
    "1110011101110111",
    "1110100000101011",
    "1110101100111111",
    "1110111011100001",
    "1111000110010110",
    "1111001010010011",
    "1111001000011101",
    "1111000100001000",
    "1110111111111101",
    "1110111110001100",
    "1110111111010100",
    "1111000010110011",
    "1111001001000010",
    "1111010011001101",
    "1111100010100010",
    "1111110111101101",
    "1111101110100101",
    "1111010011111000",
    "1110111100111000",
    "1110101110101110",
    "1110101100010100",
    "1110110100101110",
    "1111000011110011",
    "1111010011111011",
    "1111100000000111",
    "1111100101100000",
    "1111100011011100",
    "1111011011001111",
    "1111001111011010",
    "1111000011001101",
    "1110111011000100",
    "1110111011100000",
    "1111000110101100",
    "1111011011111010",
    "1111110111001111",
    "1111101101000100",
    "1111010110100111",
    "1111001001101111",
    "1111000111101000",
    "1111001110100011",
    "1111011100101000",
    "1111110000001011",
    "1111111000111001",
    "1111100000101011",
    "1111001010000110",
    "1110111000100111",
    "1110101111001111",
    "1110110000001010",
    "1110111011100110",
    "1111010000011010",
    "1111101100010111",
    "1111110100101011",
    "1111010111101101",
    "1111000001010101",
    "1110110101000011",
    "1110110011011100",
    "1110111010101101",
    "1111000111001000",
    "1111010011110110",
    "1111011101000010",
    "1111100001000011",
    "1111100000101100",
    "1111011110100001",
    "1111011101010100",
    "1111011111100011",
    "1111100110010110",
    "1111110000111101",
    "1111111101000111",
    "1111110111110011",
    "1111101111111101",
    "1111101011111000",
    "1111101010100111",
    "1111101011000011",
    "1111101101010001",
    "1111110010011111",
    "1111111100001101",
    "1111110100100110",
    "1111100000101011",
    "1111001010101000",
    "1110110110111110",
    "1110101010101010",
    "1110101001000100",
    "1110110010101100",
    "1111000100111100",
    "1111011011100000",
    "1111110010011000",
    "1111111000110111",
    "1111100111000001",
    "1111010111111010",
    "1111001011100000",
    "1111000010001111",
    "1110111101000111",
    "1110111101000101",
    "1111000010000011",
    "1111001010001100",
    "1111010011000101",
    "1111011010100110",
    "1111100000000010",
    "1111100011101001",
    "1111100101111011",
    "1111100110011001",
    "1111100011001010",
    "1111011001111100",
    "1111001010001011",
    "1110110101111011",
    "1110100001100001",
    "1110010010000000",
    "1110001011001001",
    "1110001101110000",
    "1110010111100111",
    "1110100011111011",
    "1110101111000100",
    "1110111010001110",
    "1111001001110010",
    "1111100001010101",
    "1111111110100010",
    "1111011010001011",
    "1110111000110010",
    "1110100010000011",
    "1110011011100000",
    "1110100101001011",
    "1110111001011101",
    "1111010000011110",
    "1111100101010010",
    "1111111000110111",
    "1111110000111010",
    "1111010101011000",
    "1110110101010101",
    "1110010101100111",
    "1101111101100000",
    "1101110011100010",
    "1101111010000001",
    "1110001100101110",
    "1110100011010111",
    "1110110101011010",
    "1110111101010010",
    "1110111010111000",
    "1110110001110001",
    "1110100110111001",
    "1110011110010111",
    "1110011010111000",
    "1110011111101011",
    "1110101111001100",
    "1111001001000010",
    "1111101010011000",
    "1111110010010110",
    "1111010011011101",
    "1110111110101011",
    "1110111000001011",
    "1110111111001101",
    "1111001110000111",
    "1111011101101110",
    "1111100111110111",
    "1111101010011001",
    "1111101001011110",
    "1111101011100110",
    "1111110101111101",
    "1111110110001000",
    "1111011101010010",
    "1111000111001011",
    "1110111010111100",
    "1110111100111000",
    "1111001011101000",
    "1111100001010000",
    "1111110111011111",
    "1111110110010010",
    "1111101010000010",
    "1111100011001101",
    "1111100000110001",
    "1111100001100100",
    "1111100101000101",
    "1111101100101010",
    "1111111001110100",
    "1111110011010010",
    "1111011100100001",
    "1111000101110111",
    "1110110100001000",
    "1110101010110000",
    "1110101010100110",
    "1110110010000010",
    "1110111110001010",
    "1111001011111111",
    "1111011001011000",
    "1111100101011011",
    "1111110000000110",
    "1111111010011101",
    "1111111000010001",
    "1111100100111110",
    "1111001010100101",
    "1110101010111010",
    "1110001011001110",
    "1101110001111101",
    "1101100100110001",
    "1101100111100010",
    "1101111001111100",
    "1110010111101000",
    "1110111010011001",
    "1111011011001111",
    "1111110100000010",
    "1111111111010101",
    "1111111111100110",
    "1111110011010101",
    "1111100000111110",
    "1111001101110011",
    "1110111101110111",
    "1110110011010000",
    "1110101101111011",
    "1110101101100011",
    "1110110011100001",
    "1111000001100110",
    "1111010111111100",
    "1111110100011111",
    "1111101101000111",
    "1111010010000011",
    "1110111111001101",
    "1110110111111010",
    "1110111011100101",
    "1111000110000011",
    "1111010001111110",
    "1111011010100011",
    "1111011101110000",
    "1111011100001111",
    "1111011000011000",
    "1111010101011101",
    "1111010110011011",
    "1111011110100100",
    "1111110000011100",
    "1111110011111001",
    "1111010001010101",
    "1110101101010010",
    "1110001110101000",
    "1101111011100001",
    "1101111000011000",
    "1110000101001001",
    "1110011101001010",
    "1110111011111010",
    "1111011110100110",
    "1111111101000000",
    "1111011001000001",
    "1110111000111111",
    "1110100001110000",
    "1110010110110110",
    "1110011010100101",
    "1110101011101111",
    "1111000101001000",
    "1111100010111110",
    "1111111101010111",
    "1111011110011001",
    "1111000001011111",
    "1110101000101111",
    "1110010110011000",
    "1110001011101101",
    "1110001001111010",
    "1110001111100011",
    "1110011000010101",
    "1110100000100011",
    "1110100101011011",
    "1110101000000100",
    "1110101110001100",
    "1110111100110010",
    "1111010101110110",
    "1111110111000001",
    "1111100111011001",
    "1111001110011001",
    "1111000100100100",
    "1111001100000111",
    "1111100000100111",
    "1111111001110111",
    "1111101111111111",
    "1111100010011001",
    "1111011110100100",
    "1111100011000000",
    "1111101101001100",
    "1111111010001100",
    "1111110111110101",
    "1111101001010010",
    "1111011010100101",
    "1111001100100000",
    "1111000000001111",
    "1110110111110010",
    "1110110100011101",
    "1110110101100100",
    "1110111000010101",
    "1110111001100101",
    "1110110111010101",
    "1110110001110000",
    "1110101010100110",
    "1110100100100100",
    "1110100010000101",
    "1110100011111100",
    "1110101001110100",
    "1110110010110001",
    "1110111101111101",
    "1111001100000001",
    "1111011111110001",
    "1111111011111001",
    "1111011111101001",
    "1110110110101100",
    "1110010000000101",
    "1101110011001000",
    "1101100101000000",
    "1101100111010011",
    "1101110110010110",
    "1110001011001100",
    "1110011111001000",
    "1110101101100011",
    "1110110101001101",
    "1110110111001000",
    "1110110101100100",
    "1110110011001011",
    "1110110010111101",
    "1110111000101100",
    "1111000111101111",
    "1111100000100100",
    "1111111111101010",
    "1111011110110011",
    "1111000011010111",
    "1110110010101100",
    "1110110000001000",
    "1110111010101101",
    "1111001101000100",
    "1111100000100110",
    "1111101111101111",
    "1111110111111010",
    "1111111001101001",
    "1111110111000110",
    "1111110011001001",
    "1111110000001111",
    "1111101111000101",
    "1111101111000011",
    "1111110000010010",
    "1111110101011110",
    "1111111101111001",
    "1111101000000100",
    "1111001010011000",
    "1110101010000100",
    "1110001110000000",
    "1101111100000111",
    "1101110111110100",
    "1101111111111010",
    "1110001111010010",
    "1110011111110001",
    "1110101100000101",
    "1110110010001010",
    "1110110011000001",
    "1110110010111110",
    "1110111000101010",
    "1111001000110101",
    "1111100011110110",
    "1111111001101111",
    "1111010110010110",
    "1110111000100000",
    "1110100100111011",
    "1110011101001111",
    "1110011111000101",
    "1110100110100111",
    "1110110000011100",
    "1110111001111100",
    "1111000001111101",
    "1111001000101100",
    "1111010000101001",
    "1111011110010001",
    "1111110011111111",
    "1111101111011001",
    "1111010000100111",
    "1110110110010110",
    "1110100110010011",
    "1110100011010111",
    "1110101100010100",
    "1110111011110111",
    "1111001011010100",
    "1111010100111011",
    "1111010111000001",
    "1111010110001011",
    "1111011000111111",
    "1111100100011100",
    "1111111001011000",
    "1111101100011111",
    "1111010100101111",
    "1111001000101100",
    "1111010000000011",
    "1111101011001001",
    "1111101101000000",
    "1111000011011100",
    "1110100011000011",
    "1110010010011100",
    "1110010010111110",
    "1110100011000110",
    "1110111111101100",
    "1111100101000011",
    "1111110000011011",
    "1111000100110001",
    "1110011100100001",
    "1101111100010111",
    "1101101001000010",
    "1101100101100101",
    "1101110000111011",
    "1110000110000001",
    "1110011110011011",
    "1110110100010000",
    "1111000100010011",
    "1111001110001010",
    "1111010011000000",
    "1111010101110110",
    "1111011001110010",
    "1111100000001101",
    "1111101001000011",
    "1111110010101110",
    "1111111011001100",
    "1111111110111101",
    "1111111101000000",
    "1111111110001000",
    "1111111110111011",
    "1111111100000101",
    "1111110011101000",
    "1111100110000011",
    "1111010110111110",
    "1111001010101010",
    "1111000100100100",
    "1111000110011010",
    "1111001110011100",
    "1111011000110000",
    "1111100001100110",
    "1111100110001101",
    "1111100111011110",
    "1111101010011001",
    "1111110100010001",
    "1111110111100011",
    "1111011001110100",
    "1110110111101111",
    "1110011000010001",
    "1110000010001011",
    "1101111010011110",
    "1110000001010000",
    "1110010010000011",
    "1110100110101101",
    "1110111001011001",
    "1111000110110111",
    "1111001110100011",
    "1111010001010111",
    "1111010010101110",
    "1111011000001011",
    "1111100101111100",
    "1111111101011010",
    "1111100011100111",
    "1111000010101111",
    "1110100110000011",
    "1110010010011111",
    "1110001010110111",
    "1110001110101011",
    "1110011010101101",
    "1110101010011110",
    "1110111001101000",
    "1111000101100100",
    "1111001101101101",
    "1111010010110001",
    "1111010101111001",
    "1111010111111010",
    "1111011000101010",
    "1111010111001001",
    "1111010100001011",
    "1111010011100001",
    "1111011001111001",
    "1111101010100101",
    "1111111010100001",
    "1111011001111111",
    "1110111010100101",
    "1110100011000000",
    "1110010111101010",
    "1110011000100011",
    "1110100010000110",
    "1110101111010100",
    "1110111011010001",
    "1111000011001101",
    "1111000111001000",
    "1111001000011011",
    "1111001010010001",
    "1111010000111000",
    "1111011110111010",
    "1111110100101001",
    "1111110000011011",
    "1111010101001011",
    "1110111110011011",
    "1110101111101001",
    "1110101010110101",
    "1110101111001100",
    "1110111001011011",
    "1111000101011111",
    "1111001111011010",
    "1111010101001101",
    "1111010111100000",
    "1111011000101101",
    "1111011100011110",
    "1111100101100000",
    "1111110011100100",
    "1111111100000011",
    "1111101101100100",
    "1111100100110011",
    "1111100011100010",
    "1111101000100101",
    "1111110000011011",
    "1111110110110110",
    "1111111000100110",
    "1111110100001011",
    "1111101001101000",
    "1111011001111100",
    "1111000110111110",
    "1110110011011000",
    "1110100010001011",
    "1110010110000011",
    "1110010000111101",
    "1110010011101010",
    "1110011110111011",
    "1110110100011010",
    "1111010100000000",
    "1111111010111101",
    "1111011011111100",
    "1110110111100000",
    "1110011101011011",
    "1110010001000010",
    "1110010010100010",
    "1110011101110000",
    "1110101100101101",
    "1110111010001001",
    "1111000100001011",
    "1111001110010100",
    "1111011101110111",
    "1111110101100101",
    "1111101011010111",
    "1111001010011110",
    "1110101111101001",
    "1110100001100001",
    "1110100010101111",
    "1110101111101001",
    "1110111111010010",
    "1111001000100101",
    "1111000110001110",
    "1110111001000100",
    "1110100110110100",
    "1110010110001101",
    "1110001100101110",
    "1110001100110111",
    "1110010101010011",
    "1110100100001101",
    "1110111000111010",
    "1111010010100100",
    "1111101111110100",
    "1111110001101000",
    "1111010101110110",
    "1111000001000000",
    "1110110110010010",
    "1110110101110110",
    "1110111011101011",
    "1111000011000101",
    "1111001010100101",
    "1111010011010010",
    "1111011111110000",
    "1111110001100110",
    "1111111000000100",
    "1111100000010111",
    "1111001100001001",
    "1111000001000010",
    "1111000001110100",
    "1111001101101101",
    "1111100001001111",
    "1111110111000111",
    "1111110101101000",
    "1111101000010100",
    "1111100010100001",
    "1111100100000000",
    "1111101011011001",
    "1111110111100111",
    "1111111000000001",
    "1111100011111110",
    "1111001100111010",
    "1110110101000110",
    "1110011111111101",
    "1110010001000011",
    "1110001010100011",
    "1110001100101010",
    "1110010101110110",
    "1110100011011010",
    "1110110010000110",
    "1110111111000000",
    "1111001000111110",
    "1111010000100001",
    "1111010111001101",
    "1111100000001100",
    "1111101111011100",
    "1111111000111011",
    "1111011001111101",
    "1110110111111100",
    "1110011001100011",
    "1110000100110011",
    "1101111101100000",
    "1110000100001110",
    "1110010101001011",
    "1110101010011110",
    "1110111110011111",
    "1111001101011100",
    "1111010111100101",
    "1111100000111110",
    "1111101110011101",
    "1111111101000101",
    "1111100010111000",
    "1111001000001001",
    "1110110011001101",
    "1110101001001011",
    "1110101100011110",
    "1110111011001100",
    "1111010000100011",
    "1111100111100000",
    "1111111100000110",
    "1111110011010110",
    "1111100111000111",
    "1111011111010100",
    "1111011100001111",
    "1111011110100100",
    "1111100110111010",
    "1111110100101011",
    "1111111001101101",
    "1111100110111110",
    "1111010110110100",
    "1111001100110101",
    "1111001010111010",
    "1111010000100011",
    "1111011011010001",
    "1111101000001000",
    "1111110100100110",
    "1111111110110100",
    "1111111010001010",
    "1111110110101111",
    "1111110110101000",
    "1111111000110111",
    "1111111011010101",
    "1111111011110001",
    "1111111001001000",
    "1111110100100111",
    "1111110001101010",
    "1111110100001100",
    "1111111110010001",
    "1111110000110011",
    "1111011100110000",
    "1111001011000100",
    "1111000000010010",
    "1110111110110101",
    "1111001000000100",
    "1111011011111100",
    "1111111000001000",
    "1111100111001110",
    "1111000111010110",
    "1110101100111111",
    "1110011011000010",
    "1110010011000101",
    "1110010100000000",
    "1110011001111100",
    "1110100000110000",
    "1110100110110111",
    "1110101110110001",
    "1110111100000100",
    "1111010000001111",
    "1111101001100110",
    "1111111100010011",
    "1111100111001100",
    "1111011100001100",
    "1111011101100000",
    "1111101000011111",
    "1111111000000110",
    "1111111000100001",
    "1111101100100011",
    "1111100100001110",
    "1111011110001010",
    "1111011001010110",
    "1111010101010000",
    "1111010010100001",
    "1111010010001111",
    "1111010100010000",
    "1111010111010011",
    "1111011001011101",
    "1111011000110100",
    "1111010100101010",
    "1111001110001100",
    "1111001000011110",
    "1111000111111110",
    "1111010000110011",
    "1111100100010011",
    "1111111111111101",
    "1111100010000010",
    "1111001001001011",
    "1110111011100011",
    "1110111011110111",
    "1111001000110000",
    "1111011101010001",
    "1111110010110001",
    "1111111100000111",
    "1111110010101111",
    "1111110000110001",
    "1111110001011101",
    "1111101110110100",
    "1111100100101001",
    "1111010001111110",
    "1110111001111100",
    "1110100001110110",
    "1110001111001111",
    "1110000110101100",
    "1110001001001110",
    "1110010100000001",
    "1110100010100110",
    "1110101111111101",
    "1110111000101010",
    "1110111011110111",
    "1110111011000001",
    "1110111010110010",
    "1111000000111001",
    "1111001111111011",
    "1111100110011110",
    "1111111111011000",
    "1111101100011010",
    "1111100010001111",
    "1111100011101001",
    "1111101101111011",
    "1111111011001000",
    "1111111010101111",
    "1111110111101011",
    "1111111100100001",
    "1111111000111100",
    "1111101100101010",
    "1111100010001010",
    "1111011011100011",
    "1111011000101000",
    "1111010111010110",
    "1111010101011000",
    "1111010000111001",
    "1111001001011101",
    "1110111111111010",
    "1110110101111001",
    "1110101101000000",
    "1110100110111011",
    "1110100110100010",
    "1110101111000101",
    "1111000010000011",
    "1111011110000100",
    "1111111111000110",
    "1111100000000111",
    "1111000100100101",
    "1110110001110000",
    "1110101000100000",
    "1110100111000011",
    "1110101010010100",
    "1110101111011001",
    "1110110100011101",
    "1110111001000010",
    "1110111101001110",
    "1111000001001100",
    "1111000100111100",
    "1111000111101000",
    "1111001000000110",
    "1111000101110100",
    "1111000001000111",
    "1110111011001100",
    "1110110101101100",
    "1110110001110000",
    "1110101111100110",
    "1110101110101101",
    "1110101111011010",
    "1110110100011000",
    "1111000001001000",
    "1111010111001001",
    "1111110100111101",
    "1111101001101010",
    "1111001010011001",
    "1110110010011101",
    "1110100101011000",
    "1110100011010010",
    "1110101000101101",
    "1110110000111011",
    "1110111000000100",
    "1110111100001111",
    "1110111101100110",
    "1110111101011001",
    "1110111101000000",
    "1110111110101001",
    "1111000101110100",
    "1111010100101111",
    "1111101011011101",
    "1111111000100111",
    "1111011100101110",
    "1111000110001110",
    "1110111001011000",
    "1110111000011110",
    "1111000001001101",
    "1111001111011111",
    "1111100001111101",
    "1111111000001011",
    "1111101101101110",
    "1111010000111101",
    "1110110110000000",
    "1110100001110000",
    "1110011000010011",
    "1110011100010011",
    "1110101011100000",
    "1111000000001111",
    "1111010100100101",
    "1111100100000011",
    "1111101110000101",
    "1111110101011011",
    "1111111101100001",
    "1111110110111111",
    "1111101000001110",
    "1111011000110111",
    "1111001100011011",
    "1111000101101111",
    "1111000110000000",
    "1111001011111101",
    "1111010101000011",
    "1111011110110101",
    "1111100111111011",
    "1111110000000000",
    "1111110110111011",
    "1111111100000011",
    "1111111110110000",
    "1111111110101001",
    "1111111011100110",
    "1111111000000110",
    "1111111000111010",
    "1111111110011101",
    "1111101101001100",
    "1111010101111110",
    "1110111110111011",
    "1110101110011011",
    "1110101001001110",
    "1110110000000111",
    "1110111110011110",
    "1111001101101101",
    "1111011000100101",
    "1111011101001100",
    "1111011101111011",
    "1111011111000101",
    "1111100100000000",
    "1111101110000100",
    "1111111011101000",
    "1111110111000001",
    "1111101101011100",
    "1111101001110010",
    "1111101011111011",
    "1111110010100101",
    "1111111101000011",
    "1111110100100010",
    "1111100010100111",
    "1111001111000100",
    "1110111101000111",
    "1110110000001000",
    "1110101010011110",
    "1110101100111000",
    "1110110101110100",
    "1111000001111011",
    "1111001101101101",
    "1111010110110001",
    "1111011100001100",
    "1111011110011111",
    "1111011110101001",
    "1111011101111011",
    "1111011101000010",
    "1111011100000111",
    "1111011100111111",
    "1111100010110001",
    "1111101111100001",
    "1111111100101010",
    "1111100100110111",
    "1111001110011110",
    "1110111110110110",
    "1110111010001001",
    "1111000000110101",
    "1111001110101101",
    "1111011101110101",
    "1111101001001010",
    "1111101101101010",
    "1111101101001011",
    "1111101101101001",
    "1111110100111111",
    "1111111001011001",
    "1111011111001100",
    "1111000010111101",
    "1110101100011110",
    "1110100010000011",
    "1110100101110001",
    "1110110011011101",
    "1111000011110100",
    "1111010000001100",
    "1111010101000001",
    "1111010010111000",
    "1111001100111100",
    "1111000110100100",
    "1111000010100010",
    "1111000011100110",
    "1111001100100011",
    "1111011110111111",
    "1111111001100101",
    "1111100111110101",
    "1111001011011101",
    "1110110111010011",
    "1110101111110001",
    "1110110110000001",
    "1111000110001110",
    "1111011001011000",
    "1111101010001110",
    "1111110111110101",
    "1111111011010001",
    "1111101011110011",
    "1111011000100111",
    "1111000011110011",
    "1110110010001101",
    "1110101001101010",
    "1110101110100100",
    "1111000010101100",
    "1111100100010010",
    "1111110010001110",
    "1111001000101000",
    "1110100110000011",
    "1110001111000111",
    "1110000101110010",
    "1110001001010011",
    "1110010110000000",
    "1110100110011111",
    "1110110111001001",
    "1111001000111111",
    "1111011111011111",
    "1111111100110001",
    "1111100000100001",
    "1110111101011001",
    "1110100000010101",
    "1110010000100100",
    "1110010100100100",
    "1110101101011100",
    "1111010101111100",
    "1111111011100010",
    "1111010010010000",
    "1110110110110110",
    "1110101101000010",
    "1110110100100101",
    "1111001001001100",
    "1111100011110011",
    "1111111101101100",
    "1111101110000111",
    "1111100001110000",
    "1111011100010011",
    "1111011100001001",
    "1111100000101011",
    "1111101010001101",
    "1111111000111010",
    "1111110100101010",
    "1111100001100110",
    "1111010001011010",
    "1111000111101101",
    "1111000111010110",
    "1111010000010001",
    "1111011110101001",
    "1111101101011010",
    "1111111000011001",
    "1111111110001011",
    "1111111111011111",
    "1111111101110110",
    "1111111011010001",
    "1111111010010000",
    "1111111100100101",
    "1111111100111110",
    "1111110010101001",
    "1111100101010000",
    "1111010110100000",
    "1111001000111111",
    "1110111111101001",
    "1110111100101011",
    "1111000000111110",
    "1111001011010011",
    "1111011001000110",
    "1111101000101000",
    "1111111001010100",
    "1111110100111011",
    "1111100010110011",
    "1111010010001011",
    "1111000101110100",
    "1110111111110101",
    "1111000001000011",
    "1111001000010101",
    "1111010010011001",
    "1111011011110000",
    "1111100010101110",
    "1111100111110101",
    "1111101101000010",
    "1111110011110000",
    "1111111011111011",
    "1111111011100010",
    "1111110100011010",
    "1111110000011111",
    "1111110001000000",
    "1111110110001101",
    "1111111111011110",
    "1111110100100011",
    "1111100111011000",
    "1111011010011001",
    "1111001111001000",
    "1111000110111111",
    "1111000011000101",
    "1111000011101110",
    "1111001000100011",
    "1111010000111000",
    "1111011011110111",
    "1111101000110001",
    "1111110110100110",
    "1111111100010111",
    "1111110010100001",
    "1111101110010111",
    "1111110010001011",
    "1111111111000100",
    "1111101011100110",
    "1111010000101001",
    "1110110100100101",
    "1110011100110101",
    "1110001110011110",
    "1110001101100001",
    "1110011011110000",
    "1110110111010110",
    "1111011010111100",
    "1111111111010001",
    "1111100010001111",
    "1111001101111011",
    "1111000100101100",
    "1111000100010111",
    "1111001000110000",
    "1111001101011011",
    "1111001111000100",
    "1111001100010011",
    "1111000101011101",
    "1110111011110010",
    "1110110000110101",
    "1110100110001110",
    "1110011101011001",
    "1110010111011111",
    "1110010101001110",
    "1110010110111100",
    "1110011100001111",
    "1110100011111110",
    "1110101100100110",
    "1110110100100010",
    "1110111010100101",
    "1110111110011111",
    "1111000010011101",
    "1111001011010011",
    "1111011101000100",
    "1111111000110011",
    "1111100100001110",
    "1111000000011001",
    "1110100010011100",
    "1110001111110000",
    "1110001010011101",
    "1110001111100100",
    "1110011001010001",
    "1110100010000101",
    "1110100110111001",
    "1110101000000001",
    "1110101001000110",
    "1110110000011001",
    "1111000011011111",
    "1111100011010000",
    "1111110100101011",
    "1111001100010111",
    "1110101011111101",
    "1110011001001100",
    "1110010101111110",
    "1110011110111011",
    "1110101101011100",
    "1110111011011110",
    "1111000101000011",
    "1111001000111100",
    "1111001000100011",
    "1111000110010011",
    "1111000100110100",
    "1111000110000000",
    "1111001001111001",
    "1111001111100110",
    "1111010101101100",
    "1111011011011001",
    "1111100010111110",
    "1111110000010011",
    "1111111010011011",
    "1111011110001101",
    "1110111111100011",
    "1110100100010101",
    "1110010001010010",
    "1110001001010000",
    "1110001011100001",
    "1110010011110100",
    "1110011101001100",
    "1110100011011010",
    "1110100100100100",
    "1110100001100110",
    "1110011100110111",
    "1110011001001110",
    "1110011001011101",
    "1110011110011100",
    "1110101000100010",
    "1110111000101000",
    "1111001111011111",
    "1111101100110010",
    "1111110001110100",
    "1111010001000000",
    "1110110101111110",
    "1110100100110011",
    "1110011111001010",
    "1110100011100001",
    "1110101101111111",
    "1110111010100101",
    "1111000110001101",
    "1111001111011100",
    "1111010110011101",
    "1111011011011000",
    "1111011110011001",
    "1111100000010111",
    "1111100011100001",
    "1111101010111111",
    "1111111001001101",
    "1111110000111010",
    "1111010101000011",
    "1110110111001011",
    "1110011100011100",
    "1110001010000100",
    "1110000011000011",
    "1110000110101100",
    "1110010001011010",
    "1110011110010111",
    "1110101001011101",
    "1110110000110000",
    "1110110100110110",
    "1110111001101010",
    "1111000100101010",
    "1111011001000010",
    "1111110101110011",
    "1111101001011111",
    "1111001011000100",
    "1110110100001110",
    "1110100111111001",
    "1110100101101001",
    "1110101001110111",
    "1110110001001000",
    "1110111001110100",
    "1111000100000110",
    "1111010001010101",
    "1111100010000010",
    "1111110100100000",
    "1111111010000101",
    "1111101101100010",
    "1111101001011011",
    "1111101111010001",
    "1111111110011101",
    "1111101011100111",
    "1111010011100111",
    "1110111110101110",
    "1110110001001111",
    "1110101101011011",
    "1110110011010101",
    "1111000001010000",
    "1111010101100010",
    "1111101110111111",
    "1111110011110011",
    "1111010101000011",
    "1110110111101000",
    "1110011110110101",
    "1110001101100110",
    "1110000110001110",
    "1110001001101111",
    "1110011000010011",
    "1110110001011111",
    "1111010011110001",
    "1111111100001110",
    "1111011001011110",
    "1110110010110011",
    "1110010100101100",
    "1110000010011001",
    "1101111100010111",
    "1101111111111101",
    "1110001000110000",
    "1110010010100110",
    "1110011010010110",
    "1110100000001101",
    "1110101000110010",
    "1110111010001001",
    "1111010111100111",
    "1111111111100110",
    "1111010100110011",
    "1110101110100110",
    "1110010101000000",
    "1110001011110010",
    "1110010000111110",
    "1110011101111011",
    "1110101011111100",
    "1110110110101100",
    "1110111101010110",
    "1111000000111110",
    "1111000010000101",
    "1111000000110101",
    "1110111101011011",
    "1110110111100000",
    "1110101111011001",
    "1110100110001110",
    "1110011110000000",
    "1110011001001110",
    "1110011001100101",
    "1110011111001010",
    "1110101000011011",
    "1110110011001011",
    "1110111101110000",
    "1111000111101100",
    "1111010001000101",
    "1111011010010100",
    "1111100011011000",
    "1111101011110110",
    "1111110010110011",
    "1111110111111011",
    "1111111101011111",
    "1111111000011011",
    "1111100111001000",
    "1111001110101001",
    "1110110010101100",
    "1110011001101000",
    "1110001001011101",
    "1110000110010101",
    "1110010000011110",
    "1110100011010111",
    "1110111000100101",
    "1111001001111001",
    "1111010011101001",
    "1111010101110100",
    "1111010011000101",
    "1111010000101001",
    "1111010100011000",
    "1111100000111101",
    "1111110101011010",
    "1111110010000101",
    "1111011010111111",
    "1111001001101111",
    "1111000000111011",
    "1111000000011111",
    "1111000101111100",
    "1111001110100100",
    "1111011000011101",
    "1111100011011101",
    "1111110001011111",
    "1111111011100010",
    "1111100011100100",
    "1111001001001001",
    "1110110001011001",
    "1110100001111011",
    "1110011110001111",
    "1110100110011010",
    "1110110111000100",
    "1111001011000010",
    "1111011101110011",
    "1111101101001000",
    "1111111001011010",
    "1111111011110010",
    "1111110001011011",
    "1111100111001111",
    "1111011101111010",
    "1111010110011010",
    "1111010001101001",
    "1111010000000010",
    "1111010001110100",
    "1111010110101000",
    "1111011101001111",
    "1111100011111001",
    "1111101000111110",
    "1111101011010111",
    "1111101010111001",
    "1111101000000100",
    "1111100100000000",
    "1111100000010100",
    "1111011110011011",
    "1111011111010110",
    "1111100011011010",
    "1111101010001110",
    "1111110011011110",
    "1111111111001110",
    "1111110010000000",
    "1111011111110110",
    "1111001010011000",
    "1110110010010000",
    "1110011000110101",
    "1110000000011111",
    "1101101100001010",
    "1101011110100011",
    "1101011001001011",
    "1101011011111101",
    "1101100101001101",
    "1101110010001111",
    "1101111111111111",
    "1110001101100110",
    "1110011101011110",
    "1110110010101100",
    "1111001110100011",
    "1111101110111011",
    "1111110001100011",
    "1111011001100101",
    "1111001111000101",
    "1111010101010101",
    "1111101010110010",
    "1111110110001000",
    "1111010101001101",
    "1110111001111010",
    "1110101001001001",
    "1110100100010111",
    "1110101001110100",
    "1110110101001000",
    "1111000001100001",
    "1111001011001001",
    "1111010000011010",
    "1111010100011010",
    "1111011101000000",
    "1111101110001001",
    "1111111000000011",
    "1111011010010001",
    "1110111111110110",
    "1110101111101000",
    "1110101101111111",
    "1110111010101010",
    "1111001111100100",
    "1111100100111011",
    "1111110110010110",
    "1111111010100011",
    "1111101001010001",
    "1111010010011010",
    "1110110110101000",
    "1110011010110000",
    "1110000101101100",
    "1101111110001010",
    "1110000111001001",
    "1110011101100100",
    "1110111010011110",
    "1111010101111110",
    "1111101010001100",
    "1111110101011111",
    "1111111001100101",
    "1111111001010110",
    "1111110111110011",
    "1111110111101100",
    "1111111100001000",
    "1111111000110001",
    "1111100111001101",
    "1111010001011010",
    "1110111011100000",
    "1110101010000110",
    "1110100001010101",
    "1110100100000001",
    "1110110001001000",
    "1111000100000011",
    "1111010110111111",
    "1111100101001000",
    "1111101100010111",
    "1111101110010000",
    "1111101111111001",
    "1111110111100111",
    "1111110111000111",
    "1111011110000010",
    "1111000011010000",
    "1110101110110001",
    "1110100110101111",
    "1110101100110111",
    "1110111101001010",
    "1111010000010111",
    "1111011111110000",
    "1111100111110100",
    "1111101001000101",
    "1111100111100100",
    "1111101000010111",
    "1111101111110000",
    "1111111111010101",
    "1111101011001001",
    "1111010100000101",
    "1110111111101100",
    "1110110000111101",
    "1110101000101101",
    "1110100110011010",
    "1110101000011010",
    "1110101100101011",
    "1110110001001101",
    "1110110100011000",
    "1110110100110001",
    "1110110001010100",
    "1110101010001011",
    "1110100000111001",
    "1110011000011101",
    "1110010100100111",
    "1110011000111010",
    "1110100111001011",
    "1110111110101101",
    "1111011100001001",
    "1111111010001111",
    "1111101100100011",
    "1111011100011100",
    "1111010110100101",
    "1111011000101101",
    "1111011110010111",
    "1111100011000001",
    "1111100011110001",
    "1111011111111010",
    "1111011000100101",
    "1111010000010001",
    "1111001010101111",
    "1111001100101101",
    "1111011001011000",
    "1111110000100111",
    "1111110000101011",
    "1111010000000111",
    "1110110011100010",
    "1110011111100100",
    "1110010110100101",
    "1110010111011101",
    "1110011110110110",
    "1110101001010000",
    "1110110100101001",
    "1111000001100001",
    "1111010001011111",
    "1111100101000011",
    "1111111010111000",
    "1111110000100010",
    "1111100010010101",
    "1111011111001111",
    "1111101001111111",
    "1111111101111110",
    "1111011101010100",
    "1110111011010011",
    "1110011111010010",
    "1110001110101101",
    "1110001011110101",
    "1110010110000110",
    "1110101100000010",
    "1111001011100000",
    "1111110001000011",
    "1111100111011011",
    "1111000010011101",
    "1110100100010101",
    "1110010000010100",
    "1110001000010110",
    "1110001011110101",
    "1110010111001001",
    "1110100101110001",
    "1110110100001000",
    "1111000000001111",
    "1111001010001001",
    "1111010010101100",
    "1111011011010110",
    "1111101000001000",
    "1111111101001001",
    "1111100100100010",
    "1110111111010111",
    "1110011001010001",
    "1101111001101101",
    "1101100110100000",
    "1101100011010011",
    "1101101111100100",
    "1110000110001001",
    "1110100000010100",
    "1110110111101101",
    "1111001001011011",
    "1111010111011011",
    "1111100100001101",
    "1111110000101111",
    "1111111100000001",
    "1111111101010101",
    "1111111110001011",
    "1111111001100101",
    "1111101101010101",
    "1111100011101111",
    "1111100011101111",
    "1111110000011000",
    "1111111000101011",
    "1111011110010100",
    "1111001000001000",
    "1110111010111010",
    "1110110111111111",
    "1110111101011011",
    "1111000110110010",
    "1111001111100100",
    "1111010100100100",
    "1111010100100010",
    "1111010000100001",
    "1111001010110111",
    "1111000110101010",
    "1111000111011011",
    "1111001111101001",
    "1111011111110011",
    "1111110101110110",
    "1111110010001110",
    "1111011100111111",
    "1111001101101000",
    "1111000101010000",
    "1111000010101110",
    "1111000011100010",
    "1111000101100111",
    "1111000111110111",
    "1111001010100110",
    "1111001110111111",
    "1111010101011111",
    "1111011101100000",
    "1111100101000001",
    "1111101001011010",
    "1111101000110111",
    "1111100010111011",
    "1111011000110000",
    "1111001101000000",
    "1111000010111000",
    "1110111101000111",
    "1110111100110101",
    "1111000001010010",
    "1111001000010001",
    "1111010000010101",
    "1111011010101101",
    "1111101001010110",
    "1111111100110011",
    "1111101100100001",
    "1111010110001001",
    "1111000100001010",
    "1110111001111100",
    "1110111001010001",
    "1111000000110000",
    "1111001100001100",
    "1111010111010000",
    "1111011110100110",
    "1111100001001111",
    "1111100000001010",
    "1111011100111100",
    "1111011001010011",
    "1111010110101010",
    "1111010101010000",
    "1111010100100010",
    "1111010011111000",
    "1111010010101110",
    "1111010001011111",
    "1111010010100001",
    "1111011000011010",
    "1111100100000000",
    "1111110011111111",
    "1111111010111001",
    "1111101100110101",
    "1111100101011000",
    "1111100110100000",
    "1111101110111111",
    "1111111010101010",
    "1111111011011101",
    "1111110111100100",
    "1111111011010000",
    "1111111010111110",
    "1111101110111010",
    "1111100101101100",
    "1111100011111100",
    "1111101011101111",
    "1111111011111100",
    "1111101111001101",
    "1111011011001110",
    "1111001101011100",
    "1111001010000100",
    "1111010010111001",
    "1111100110101101",
    "1111111110001101",
    "1111100000111011",
    "1111000110100000",
    "1110110010111001",
    "1110101000010110",
    "1110100111001011",
    "1110101110001100",
    "1110111011001110",
    "1111001011111000",
    "1111011101101001",
    "1111101110010000",
    "1111111100011010",
    "1111110110101000",
    "1111101000010101",
    "1111010110101010",
    "1111000001010000",
    "1110101010100101",
    "1110010110111011",
    "1110001010100101",
    "1110001000011101",
    "1110010000010010",
    "1110100000011010",
    "1110111000011110",
    "1111010111100111",
    "1111111011101110",
    "1111011110100011",
    "1110111100011110",
    "1110100011000011",
    "1110010110000100",
    "1110010111001000",
    "1110100011101111",
    "1110110110101100",
    "1111001010100000",
    "1111011010110000",
    "1111100101100111",
    "1111101100001011",
    "1111110001011011",
    "1111111001001011",
    "1111111010101010",
    "1111101011101011",
    "1111011101010110",
    "1111010011011111",
    "1111010000001100",
    "1111010010011101",
    "1111010110111110",
    "1111011010000100",
    "1111011001101011",
    "1111010110000001",
    "1111010001000011",
    "1111001101001111",
    "1111001100101000",
    "1111010001011111",
    "1111011101011110",
    "1111110000010010",
    "1111111000011101",
    "1111100000111011",
    "1111001101100011",
    "1111000001110001",
    "1110111111101011",
    "1111000110101100",
    "1111010100000011",
    "1111100110001011",
    "1111111100011010",
    "1111101010010111",
    "1111001111101001",
    "1110110110001101",
    "1110100001010100",
    "1110010011011111",
    "1110001110110101",
    "1110010011001101",
    "1110011101011001",
    "1110101001010011",
    "1110110011000000",
    "1110111000000001",
    "1110111000010101",
    "1110110101100000",
    "1110110010010100",
    "1110110001001100",
    "1110110010100100",
    "1110110101100100",
    "1110111001101011",
    "1110111111110000",
    "1111001001011011",
    "1111010111111111",
    "1111101010101100",
    "1111111110000111",
    "1111110010001110",
    "1111101001111000",
    "1111101001010111",
    "1111101101110000",
    "1111110010000100",
    "1111110001110100",
    "1111101010110111",
    "1111011110010100",
    "1111001111101100",
    "1111000010111101",
    "1110111010110000",
    "1110110111011011",
    "1110110111010011",
    "1110111000001001",
    "1110111000111110",
    "1110111011000001",
    "1111000001001101",
    "1111001110010010",
    "1111100010101001",
    "1111111011000011",
    "1111101110001000",
    "1111011110011001",
    "1111011000110100",
    "1111011101000101",
    "1111101000000011",
    "1111110101001000",
    "1111111111100000",
    "1111110111111000",
    "1111110011111111",
    "1111110010101011",
    "1111110010100001",
    "1111110010100010",
    "1111110010010011",
    "1111110001101101",
    "1111110000011011",
    "1111101101101010",
    "1111101000100111",
    "1111100001010101",
    "1111011001011000",
    "1111010011110110",
    "1111010100100111",
    "1111011110001001",
    "1111110000000010",
    "1111111001000010",
    "1111100010100010",
    "1111010001101100",
    "1111001010000110",
    "1111001100100001",
    "1111010110111001",
    "1111100100111110",
    "1111110010010000",
    "1111111010111111",
    "1111111101001101",
    "1111111001010100",
    "1111110001101110",
    "1111101001111110",
    "1111100101001110",
    "1111100100111110",
    "1111101000101101",
    "1111101110010111",
    "1111110010111011",
    "1111110011100100",
    "1111101110100001",
    "1111100011100100",
    "1111010100001011",
    "1111000011100110",
    "1110110101100101",
    "1110101101111010",
    "1110110000010101",
    "1110111111101001",
    "1111011011110011",
    "1111111110100100",
    "1111010101110110",
    "1110110001000011",
    "1110010110000100",
    "1110001000001011",
    "1110000110101100",
    "1110001101100110",
    "1110010111111001",
    "1110100001100110",
    "1110101011001111",
    "1110111001011101",
    "1111010000000000",
    "1111101111111000",
    "1111101010001110",
    "1111000101100101",
    "1110101001100101",
    "1110011011100101",
    "1110011100110101",
    "1110101000110111",
    "1110111000110100",
    "1111000110001101",
    "1111001101010110",
    "1111001110100100",
    "1111001100001010",
    "1111001000110010",
    "1111001000001011",
    "1111001110001111",
    "1111011101001010",
    "1111110100101101",
    "1111101110001000",
    "1111010000101110",
    "1110111000010001",
    "1110101001000110",
    "1110100101100100",
    "1110101101000000",
    "1110111101100100",
    "1111010101000101",
    "1111110000000100",
    "1111110100111101",
    "1111011101101110",
    "1111001110000101",
    "1111001000001000",
    "1111001100100110",
    "1111011011001010",
    "1111110010010001",
    "1111110000000001",
    "1111001110011100",
    "1110101100101000",
    "1110001110110101",
    "1101111001001011",
    "1101101110010111",
    "1101101110111010",
    "1101111001001110",
    "1110001010000110",
    "1110011101100001",
    "1110110001100001",
    "1111000111000100",
    "1111100000010111",
    "1111111110001010",
    "1111100000111110",
    "1111000000111000",
    "1110100110010000",
    "1110010101011010",
    "1110010000100011",
    "1110010110100000",
    "1110100011011101",
    "1110110010110011",
    "1111000000111101",
    "1111001100011011",
    "1111010101010010",
    "1111011011110010",
    "1111100000011100",
    "1111100011100001",
    "1111100101000011",
    "1111100101011000",
    "1111100110010010",
    "1111101010010111",
    "1111110011110110",
    "1111111100101111",
    "1111101001011111",
    "1111010110011000",
    "1111000111101100",
    "1110111111110110",
    "1110111110010110",
    "1110111111111101",
    "1111000000110000",
    "1110111110010001",
    "1110111000010011",
    "1110110000111001",
    "1110101011000010",
    "1110101001000111",
    "1110101011111010",
    "1110110010000101",
    "1110111001001001",
    "1110111111000101",
    "1111000010111101",
    "1111000101001000",
    "1111001000011011",
    "1111010001010100",
    "1111100010111110",
    "1111111101010110",
    "1111100010110110",
    "1111000011000110",
    "1110101000110101",
    "1110011000100011",
    "1110010100100000",
    "1110011011101000",
    "1110101010010011",
    "1110111011111101",
    "1111001100011011",
    "1111011000110100",
    "1111100001100110",
    "1111101010101011",
    "1111111000100100",
    "1111110010011000",
    "1111010111011011",
    "1110111011001001",
    "1110100011001011",
    "1110010100110001",
    "1110010010011101",
    "1110011010010110",
    "1110100111101111",
    "1110110101100010",
    "1111000001011100",
    "1111001101101000",
    "1111011101100001",
    "1111110011000011",
    "1111110010010001",
    "1111010110101000",
    "1110111111111011",
    "1110110011010011",
    "1110110011010000",
    "1110111111011010",
    "1111010101101010",
    "1111110010000101",
    "1111110000001010",
    "1111010101100100",
    "1111000001110110",
    "1110110111101000",
    "1110110111100111",
    "1111000000010101",
    "1111001101101000",
    "1111011011111101",
    "1111101011111001",
    "1111111111111001",
    "1111100110001001",
    "1111000111011111",
    "1110101000101101",
    "1110001111010110",
    "1110000000110001",
    "1110000000111101",
    "1110001110110110",
    "1110100101011101",
    "1110111111011111",
    "1111011010000111",
    "1111110101011011",
    "1111101101000101",
    "1111001100111100",
    "1110101011101011",
    "1110001101011110",
    "1101111000010001",
    "1101110001001000",
    "1101111001011011",
    "1110001110100011",
    "1110101011000100",
    "1111001000011101",
    "1111100001101110",
    "1111110100011101",
    "1111111111100100",
    "1111111001000010",
    "1111110110010011",
    "1111110100110101",
    "1111110000100000",
    "1111100110010010",
    "1111010101111100",
    "1111000010010010",
    "1110110000010010",
    "1110100101000000",
    "1110100100011101",
    "1110101111110011",
    "1111000011010000",
    "1111010111001011",
    "1111100011100111",
    "1111100011110011",
    "1111011000001001",
    "1111000101010101",
    "1110110010000000",
    "1110100100011101",
    "1110100000000101",
    "1110100100000110",
    "1110101100101011",
    "1110110101001101",
    "1110111011001110",
    "1111000000010100",
    "1111001001011110",
    "1111011011000110",
    "1111110101111110",
    "1111101001101010",
    "1111001010111111",
    "1110110100111110",
    "1110101100011100",
    "1110110010100010",
    "1111000011100111",
    "1111011001101010",
    "1111101111010000",
    "1111111110011110",
    "1111101111001010",
    "1111100000110011",
    "1111010001111000",
    "1111000010000011",
    "1110110010110100",
    "1110100110101111",
    "1110100000000111",
    "1110011111111111",
    "1110100101011101",
    "1110101101111111",
    "1110110110110010",
    "1110111110000111",
    "1111000011010111",
    "1111000111011101",
    "1111001101111010",
    "1111011010110101",
    "1111110000010011",
    "1111110011000000",
    "1111010100000001",
    "1110111001001110",
    "1110101000001001",
    "1110100011111011",
    "1110101010111111",
    "1110110111111111",
    "1111000100110110",
    "1111001100101011",
    "1111001101010010",
    "1111000111110010",
    "1110111110101110",
    "1110110101100000",
    "1110101111001000",
    "1110101100110010",
    "1110101110011001",
    "1110110011000011",
    "1110111001000010",
    "1110111110110110",
    "1111000011100110",
    "1111000110111001",
    "1111001000101000",
    "1111001000110111",
    "1111001000000110",
    "1111000111101101",
    "1111001010010011",
    "1111010010111001",
    "1111100011100100",
    "1111111100001010",
    "1111100101110111",
    "1111000110101000",
    "1110101010101111",
    "1110010110011011",
    "1110001100010100",
    "1110001100100011",
    "1110010101010010",
    "1110100011100100",
    "1110110100100000",
    "1111000101101100",
    "1111010101010000",
    "1111100001111101",
    "1111101011001010",
    "1111110000101001",
    "1111110010110110",
    "1111110101001101",
    "1111111101001011",
    "1111110001101100",
    "1111010111100101",
    "1110111000111100",
    "1110011101010100",
    "1110001011101011",
    "1110001000011010",
    "1110010011001111",
    "1110100110100111",
    "1110111011101011",
    "1111001100111100",
    "1111010111111001",
    "1111011111001000",
    "1111101000010000",
    "1111110111101101",
    "1111110001011010",
    "1111010111011101",
    "1111000010001101",
    "1110111000011000",
    "1110111100111111",
    "1111001101100110",
    "1111100010100001",
    "1111110010011110",
    "1111110111010001",
    "1111101111110001",
    "1111100000000010",
    "1111001110110011",
    "1111000010100100",
    "1111000000011010",
    "1111001010010001",
    "1111011110011011",
    "1111111000101110",
    "1111101100011110",
    "1111010110010011",
    "1111000111101000",
    "1111000000111110",
    "1111000000110110",
    "1111000100100111",
    "1111001001101000",
    "1111001101101101",
    "1111001111100001",
    "1111001110111101",
    "1111001100111100",
    "1111001011001001",
    "1111001011111111",
    "1111010001111011",
    "1111011110111111",
    "1111110011110101",
    "1111110000110101",
    "1111010001111110",
    "1110110011011000",
    "1110011000111010",
    "1110000101101001",
    "1101111011000111",
    "1101111001000001",
    "1101111101111010",
    "1110001000111001",
    "1110011001111010",
    "1110110000010111",
    "1111001001110100",
    "1111100010001101",
    "1111110101000100",
    "1111111111000100",
    "1111111111010110",
    "1111111000001111",
    "1111101110110000",
    "1111101000101100",
    "1111101010010111",
    "1111110101001111",
    "1111111000001010",
    "1111100000111110",
    "1111001000100011",
    "1110110001110000",
    "1110011110010010",
    "1110001111010111",
    "1110000101111011",
    "1110000010010111",
    "1110000100101110",
    "1110001100001001",
    "1110010111001110",
    "1110100101100000",
    "1110110111100010",
    "1111001101110010",
    "1111100111111110",
    "1111111011011101",
    "1111011111001000",
    "1111000101101001",
    "1110110001001100",
    "1110100010100111",
    "1110011000111110",
    "1110010010100010",
    "1110001101111000",
    "1110001010010100",
    "1110001000001011",
    "1110000111110101",
    "1110001001101111",
    "1110001110001001",
    "1110010100101010",
    "1110011100011011",
    "1110100100010111",
    "1110101011100011",
    "1110110001010111",
    "1110110101101010",
    "1110111000101111",
    "1110111010111111",
    "1110111100111111",
    "1110111111101011",
    "1111000101101111",
    "1111010011100010",
    "1111101100000101",
    "1111110000110100",
    "1111000111010011",
    "1110011110101011",
    "1101111110101110",
    "1101101101011011",
    "1101101101000010",
    "1101111010101011",
    "1110010000001101",
    "1110100111000110",
    "1110111010001011",
    "1111000111101101",
    "1111010000100100",
    "1111010111101100",
    "1111100010111110",
    "1111110111010100",
    "1111101010101011",
    "1111000110001110",
    "1110100010000010",
    "1110000101100000",
    "1101110110000000",
    "1101110110000011",
    "1110000011101100",
    "1110011001110100",
    "1110110101100000",
    "1111010101111001",
    "1111111010001000",
    "1111011110110000",
    "1110111000100010",
    "1110011000001100",
    "1110000010001011",
    "1101111010010011",
    "1110000000100111",
    "1110010001000000",
    "1110100111101010",
    "1111000001110000",
    "1111011100101110",
    "1111110110110101",
    "1111110010110111",
    "1111100100001010",
    "1111011111111111",
    "1111101000101101",
    "1111111101001010",
    "1111101000101111",
    "1111010000110110",
    "1111000010001111",
    "1111000001000111",
    "1111001100110111",
    "1111100001011010",
    "1111111000111001",
    "1111110010010010",
    "1111100010111001",
    "1111011000101101",
    "1111010010001111",
    "1111001101011011",
    "1111001001000010",
    "1111000101100100",
    "1111000100001000",
    "1111000101111100",
    "1111001011001010",
    "1111010010110001",
    "1111011011001010",
    "1111100010110100",
    "1111101000101110",
    "1111101100110001",
    "1111101111111110",
    "1111110100000001",
    "1111111010100011",
    "1111111011100111",
    "1111101111000100",
    "1111100001001010",
    "1111010011111110",
    "1111001001011000",
    "1111000010001011",
    "1110111101110101",
    "1110111010100000",
    "1110110110010010",
    "1110110000001101",
    "1110101000011110",
    "1110100000011010",
    "1110011010000001",
    "1110010111000100",
    "1110011000010001",
    "1110011101010001",
    "1110100100110111",
    "1110101110100011",
    "1110111100010011",
    "1111010001000010",
    "1111101110000000",
    "1111101110011110",
    "1111001001100011",
    "1110101010000001",
    "1110010101100101",
    "1110001111011010",
    "1110010110000100",
    "1110100100000101",
    "1110110011001010",
    "1110111110101110",
    "1111000101111011",
    "1111001011000111",
    "1111010001001100",
    "1111011001110010",
    "1111100100011000",
    "1111101101111010",
    "1111110011001001",
    "1111110010100111",
    "1111101101001111",
    "1111100110001011",
    "1111100001001100",
    "1111100000011111",
    "1111100011111000",
    "1111101000110000",
    "1111101100001111",
    "1111101100101001",
    "1111101011010000",
    "1111101100110111",
    "1111110110100111",
    "1111110100111101",
    "1111010111010110",
    "1110110110001000",
    "1110011000010110",
    "1110000100010010",
    "1101111101010001",
    "1110000001110001",
    "1110001101000010",
    "1110011010001110",
    "1110100101101010",
    "1110101111000010",
    "1110111010011001",
    "1111001100010011",
    "1111100110101000",
    "1111111000110011",
    "1111011000110100",
    "1111000000111110",
    "1110110110101100",
    "1110111011111101",
    "1111001101011100",
    "1111100011101110",
    "1111110111100000",
    "1111111011110111",
    "1111110111011110",
    "1111111001000111",
    "1111111110010001",
    "1111111011010101",
    "1111110101011011",
    "1111101111111111",
    "1111101010101001",
    "1111100101011010",
    "1111100000001010",
    "1111011011011001",
    "1111010111101111",
    "1111010101001001",
    "1111010011000001",
    "1111010000010100",
    "1111001101001001",
    "1111001101100000",
    "1111010110011010",
    "1111101010010000",
    "1111111000010000",
    "1111010111000001",
    "1110111001101111",
    "1110100110101101",
    "1110100001100001",
    "1110101000101010",
    "1110110110010011",
    "1111000100001011",
    "1111001101100110",
    "1111010001001000",
    "1111010000100100",
    "1111001101111111",
    "1111001100101011",
    "1111010001110000",
    "1111011111101001",
    "1111110101010010",
    "1111110001000100",
    "1111011001101010",
    "1111001001110010",
    "1111000100110011",
    "1111001011110010",
    "1111011011101101",
    "1111101111001100",
    "1111111111000000",
    "1111110011000000",
    "1111101100000010",
    "1111100101011010",
    "1111011011000100",
    "1111001010110000",
    "1110110101110110",
    "1110100001010100",
    "1110010010010100",
    "1110001101000010",
    "1110010010101100",
    "1110011111111000",
    "1110101111001101",
    "1110111100001010",
    "1111000110011101",
    "1111010010011001",
    "1111100011111001",
    "1111111100010101",
    "1111100110000100",
    "1111001000101100",
    "1110110001111110",
    "1110100111000011",
    "1110101001110010",
    "1110110111000110",
    "1111001000110010",
    "1111011000111010",
    "1111100011101001",
    "1111101000100100",
    "1111101001001101",
    "1111100111011110",
    "1111100110100101",
    "1111101010010000",
    "1111110100100001",
    "1111111010101010",
    "1111100101111110",
    "1111010001101011",
    "1111000001101100",
    "1110111001000110",
    "1110111001101011",
    "1111000011000001",
    "1111010010101110",
    "1111100100101100",
    "1111110100011010",
    "1111111110100101",
    "1111111111000010",
    "1111111010001101",
    "1111101011011101",
    "1111010111111100",
    "1111000011110001",
    "1110110010111011",
    "1110100111110100",
    "1110100011000101",
    "1110100100100100",
    "1110101011000111",
    "1110110100110001",
    "1110111111101110",
    "1111001100101011",
    "1111011111000000",
    "1111111001001010",
    "1111100101101111",
    "1111000010000011",
    "1110100010100100",
    "1110001110110000",
    "1110001100101011",
    "1110011110011100",
    "1111000000000000",
    "1111101001000011",
    "1111101111110101",
    "1111010010101100",
    "1111000011010111",
    "1111000001001111",
    "1111001000011110",
    "1111010011011100",
    "1111011100111111",
    "1111100010001101",
    "1111100010101001",
    "1111100001010010",
    "1111100100000110",
    "1111110000001100",
    "1111111000101010",
    "1111011000011010",
    "1110110100010011",
    "1110010011101100",
    "1101111110000111",
    "1101111000110010",
    "1110000011010011",
    "1110011000111001",
    "1110110100011111",
    "1111010010100111",
    "1111110001011011",
    "1111110000100111",
    "1111010110001110",
    "1111000010001111",
    "1110110111001001",
    "1110110111010001",
    "1111000011101100",
    "1111011011000100",
    "1111111010001001",
    "1111100011010011",
    "1111000001001000",
    "1110100010001000",
    "1110001000110100",
    "1101110111011000",
    "1101101111001010",
    "1101110000000010",
    "1101111000011011",
    "1110000101101110",
    "1110010100101010",
    "1110100010100001",
    "1110101101011100",
    "1110110100111110",
    "1110111100011011",
    "1111001001100101",
    "1111011111111011",
    "1111111110101110",
    "1111011111001111",
    "1111000001101001",
    "1110101110110011",
    "1110101010111100",
    "1110110110001000",
    "1111001011010110",
    "1111100011111100",
    "1111111001110010",
    "1111110101011110",
    "1111100110101000",
    "1111010101101001",
    "1111000001001000",
    "1110101010110111",
    "1110010111111111",
    "1110001110010100",
    "1110010000111101",
    "1110011111010010",
    "1110110011110001",
    "1111000110000011",
    "1111001111011110",
    "1111001101101110",
    "1111000011101001",
    "1110110110101100",
    "1110101011101010",
    "1110100101111001",
    "1110100111110001",
    "1110110010001011",
    "1111000100100010",
    "1111011100101101",
    "1111110110111011",
    "1111110001000001",
    "1111011111010010",
    "1111010111110101",
    "1111011101001001",
    "1111101110101110",
    "1111110110111001",
    "1111011001100000",
    "1110111111010001",
    "1110101101000111",
    "1110100110010011",
    "1110101011110101",
    "1110111100001111",
    "1111010100011100",
    "1111110000011001",
    "1111110100000011",
    "1111011100100110",
    "1111001011111101",
    "1111000011100111",
    "1111000011010111",
    "1111001001001110",
    "1111010001101110",
    "1111011001001001",
    "1111011100101101",
    "1111011011010011",
    "1111010110000000",
    "1111010000001111",
    "1111001110111011",
    "1111010110001011",
    "1111100111001010",
    "1111111111100100",
    "1111100101100000",
    "1111001110001100",
    "1110111111011110",
    "1110111100010100",
    "1111000101010111",
    "1111011000111001",
    "1111110011101100",
    "1111101101110011",
    "1111001111000101",
    "1110110011100001",
    "1110011110100011",
    "1110010011110110",
    "1110010110011000",
    "1110100111010101",
    "1111000101001101",
    "1111101011110011",
    "1111101011000011",
    "1111000110100100",
    "1110101100111100",
    "1110100001011110",
    "1110100011101111",
    "1110110000010100",
    "1111000010001101",
    "1111010101101100",
    "1111101001101000",
    "1111111110011011",
    "1111101011011111",
    "1111010100111001",
    "1111000000000011",
    "1110110000001000",
    "1110101000100010",
    "1110101011011001",
    "1110111000001100",
    "1111001100010100",
    "1111100100000110",
    "1111111100010100",
    "1111101100111110",
    "1111011000101010",
    "1111000111010011",
    "1110111001001110",
    "1110101111000000",
    "1110101001011101",
    "1110101001001011",
    "1110101110011011",
    "1110111000110101",
    "1111001000101100",
    "1111011111001100",
    "1111111101000111",
    "1111011110101000",
    "1110110111110001",
    "1110010100010010",
    "1101111010101111",
    "1101110000000111",
    "1101110110001011",
    "1110001001111010",
    "1110100100111100",
    "1110111111111011",
    "1111010100101110",
    "1111100000000011",
    "1111100001111110",
    "1111011110110110",
    "1111011110001001",
    "1111100101100100",
    "1111110110011110",
    "1111110010011011",
    "1111011011111111",
    "1111001101001001",
    "1111001010100010",
    "1111010101000011",
    "1111101011010110",
    "1111110100110001",
    "1111001110111111",
    "1110101000000100",
    "1110000101101010",
    "1101101101010100",
    "1101100010111110",
    "1101101000001011",
    "1101111010101111",
    "1110010111000011",
    "1110111010101111",
    "1111100011010010",
    "1111110010001101",
    "1111001001011101",
    "1110100111011011",
    "1110010000001101",
    "1110000110000110",
    "1110001001111111",
    "1110011000111111",
    "1110101101110010",
    "1111000010110011",
    "1111010010111110",
    "1111011100000010",
    "1111011110010110",
    "1111011100001111",
    "1111011001011110",
    "1111011001101111",
    "1111100000000111",
    "1111101110110010",
    "1111111010010111",
    "1111011110001001",
    "1111000001001000",
    "1110101000100000",
    "1110011001000001",
    "1110010101110001",
    "1110011110000010",
    "1110101101011100",
    "1110111110010001",
    "1111001011011110",
    "1111010010011100",
    "1111010011000000",
    "1111001110100100",
    "1111000111011101",
    "1110111111110110",
    "1110111010001001",
    "1110111001011101",
    "1111000000100011",
    "1111010000100001",
    "1111101000000001",
    "1111111100011011",
    "1111100001011001",
    "1111001011001111",
    "1110111100111111",
    "1110110110110010",
    "1110110110100111",
    "1110111001011011",
    "1110111100100001",
    "1110111110011100",
    "1110111110111101",
    "1110111110010111",
    "1110111101001001",
    "1110111011101111",
    "1110111010101010",
    "1110111010011110",
    "1110111100100001",
    "1111000010101111",
    "1111001111011010",
    "1111100011101001",
    "1111111110011110",
    "1111100010111000",
    "1111000100010101",
    "1110101010001100",
    "1110011000000001",
    "1110001111101000",
    "1110010000101011",
    "1110011000111010",
    "1110100101001110",
    "1110110010011010",
    "1110111101101000",
    "1111000110011111",
    "1111001111011001",
    "1111011011010110",
    "1111101011111000",
    "1111111111110110",
    "1111101011001001",
    "1111011010000001",
    "1111001111111011",
    "1111001110101001",
    "1111010101000101",
    "1111100000011001",
    "1111101101011001",
    "1111111001010010",
    "1111111101101011",
    "1111111000001010",
    "1111110110010100",
    "1111110111100010",
    "1111111011001011",
    "1111111111001110",
    "1111111000100110",
    "1111110001111101",
    "1111101100011010",
    "1111101001001100",
    "1111101001000010",
    "1111101011110101",
    "1111110001000100",
    "1111111000010011",
    "1111111110000110",
    "1111110001010101",
    "1111100000110110",
    "1111001101001111",
    "1110111000010011",
    "1110100100111110",
    "1110010110101010",
    "1110010000110000",
    "1110010101101111",
    "1110100101111001",
    "1110111110110000",
    "1111011011011001",
    "1111110101110110",
    "1111110111001101",
    "1111101110111011",
    "1111110001001110",
    "1111111010110001",
    "1111111010001111",
    "1111110101000110",
    "1111111011101111",
    "1111101111101010",
    "1111001111111011",
    "1110101100001100",
    "1110001101100011",
    "1101111011110011",
    "1101111010111000",
    "1110001001010011",
    "1110100000110101",
    "1110111001110010",
    "1111001101101101",
    "1111011001100011",
    "1111011111111000",
    "1111100111010000",
    "1111110101101111",
    "1111110001111111",
    "1111010010110001",
    "1110110011100100",
    "1110011100001111",
    "1110010011011000",
    "1110011100000111",
    "1110110100000101",
    "1111010101001110",
    "1111111000001011",
    "1111101001110110",
    "1111010101000001",
    "1111001010011101",
    "1111001000101000",
    "1111001011001111",
    "1111001101010111",
    "1111001011101000",
    "1111000100110001",
    "1110111010011001",
    "1110101111101011",
    "1110100111001110",
    "1110100010011111",
    "1110100001010111",
    "1110100010101110",
    "1110100100111011",
    "1110100110011000",
    "1110100110010010",
    "1110100101000101",
    "1110100100000101",
    "1110100101010101",
    "1110101011011011",
    "1110110111111010",
    "1111001010010011",
    "1111011111111011",
    "1111110100100000",
    "1111111100001011",
    "1111110100011111",
    "1111110100000011",
    "1111110111011100",
    "1111111001100001",
    "1111110101110001",
    "1111101001101111",
    "1111010110000011",
    "1110111110000100",
    "1110100110011011",
    "1110010011011100",
    "1110000111110111",
    "1110000100011010",
    "1110001000010101",
    "1110010001110001",
    "1110011110010110",
    "1110101011111111",
    "1110111001000111",
    "1111000100100100",
    "1111001101101000",
    "1111010011110110",
    "1111010111001001",
    "1111011001110111",
    "1111100000111110",
    "1111110000011111",
    "1111110110111100",
    "1111011000111110",
    "1110111100010110",
    "1110100111111110",
    "1110100000110000",
    "1110100111110101",
    "1110111010001100",
    "1111010011110011",
    "1111110001001001",
    "1111110000101001",
    "1111010011010111",
    "1110111000101111",
    "1110100010111101",
    "1110010011111110",
    "1110001101100001",
    "1110010000010001",
    "1110011011101000",
    "1110101111000000",
    "1111001000100011",
    "1111100100110111",
    "1111111111101011",
    "1111101010111010",
    "1111011101001001",
    "1111010111100101",
    "1111011001111001",
    "1111100010010101",
    "1111101110001001",
    "1111111010100101",
    "1111111010100000",
    "1111110010100101",
    "1111101101111010",
    "1111101011100101",
    "1111101010000110",
    "1111101000001011",
    "1111100101010011",
    "1111100001110100",
    "1111011110110001",
    "1111011110000100",
    "1111100001111000",
    "1111101100011011",
    "1111111110111001",
    "1111100111101100",
    "1111001011001010",
    "1110110001001000",
    "1110011111001101",
    "1110011000110111",
    "1110011110101000",
    "1110101110100110",
    "1111000101011101",
    "1111100000001010",
    "1111111100101010",
    "1111100110011000",
    "1111001010000111",
    "1110101111110001",
    "1110011001011101",
    "1110001001111100",
    "1110000011110011",
    "1110001000000100",
    "1110010101001110",
    "1110101000101111",
    "1111000001110000",
    "1111100000001100",
    "1111111100100010",
    "1111010110001110",
    "1110110000101011",
    "1110010000100011",
    "1101111010011011",
    "1101110001010000",
    "1101110101001011",
    "1110000101100100",
    "1110100001000011",
    "1111000100011000",
    "1111101011001111",
    "1111101111101100",
    "1111010010001000",
    "1111000000010001",
    "1110111100000010",
    "1111000100000110",
    "1111010011110011",
    "1111100101100101",
    "1111110110100100",
    "1111110111111101",
    "1111100011100110",
    "1111001011100101",
    "1110110001100001",
    "1110011001110000",
    "1110001010001001",
    "1110000111110101",
    "1110010100110110",
    "1110101101100110",
    "1111001010111101",
    "1111100101011011",
    "1111111000011011",
    "1111111010010100",
    "1111101101100100",
    "1111011101010001",
    "1111001000010000",
    "1110110001100010",
    "1110011111000111",
    "1110010110100000",
    "1110011011000110",
    "1110101011111100",
    "1111000011110011",
    "1111011011111010",
    "1111101111101111",
    "1111111111101111",
    "1111101110000101",
    "1111010111101000",
    "1110111011111101",
    "1110011110011111",
    "1110000101110001",
    "1101111000010110",
    "1101111010000001",
    "1110001001011001",
    "1110100000010010",
    "1110110111001011",
    "1111001000011000",
    "1111010001110000",
    "1111010100100111",
    "1111010011010111",
    "1111010000111001",
    "1111010001001000",
    "1111011000000011",
    "1111100111101010",
    "1111111111010011",
    "1111100100011100",
    "1111001000110100",
    "1110110010110100",
    "1110100110110010",
    "1110100110110001",
    "1110110000011110",
    "1110111110011011",
    "1111001010010100",
    "1111001111011110",
    "1111001101000000",
    "1111000100111011",
    "1110111010111000",
    "1110110011010101",
    "1110110001001101",
    "1110110100111001",
    "1110111100110000",
    "1111000110000100",
    "1111001111010111",
    "1111011001011101",
    "1111100110111010",
    "1111111001111100",
    "1111101101001111",
    "1111010000111011",
    "1110110101000001",
    "1110011110010110",
    "1110010001000101",
    "1110001111000111",
    "1110010110101100",
    "1110100011010111",
    "1110110000000011",
    "1110111001000010",
    "1110111100111101",
    "1110111100100110",
    "1110111001111101",
    "1110110111110010",
    "1110111001110010",
    "1111000011110100",
    "1111010111101010",
    "1111110100000001",
    "1111101011000001",
    "1111001010111111",
    "1110110000111011",
    "1110100000100110",
    "1110011011010011",
    "1110011110111101",
    "1110100111110010",
    "1110110010101110",
    "1110111110111111",
    "1111001101110101",
    "1111100000011001",
    "1111110101110011",
    "1111110100100101",
    "1111100011000000",
    "1111011001101010",
    "1111011010111000",
    "1111100101110001",
    "1111110101111101",
    "1111111010101010",
    "1111110001001001",
    "1111101111100000",
    "1111110100101000",
    "1111111101011110",
    "1111111001001010",
    "1111110001101001",
    "1111101100101010",
    "1111101001000110",
    "1111100100100111",
    "1111011101000111",
    "1111010010001111",
    "1111000101011111",
    "1110111001100111",
    "1110110001010000",
    "1110101101111011",
    "1110101111110011",
    "1110110101110111",
    "1110111110011111",
    "1111000111111110",
    "1111010001100110",
    "1111011110000000",
    "1111110001100111",
    "1111110001110100",
    "1111001110001001",
    "1110101000111001",
    "1110001001110101",
    "1101110111011101",
    "1101110101110010",
    "1110000100001000",
    "1110011100011011",
    "1110110110111110",
    "1111001101000111",
    "1111011101010010",
    "1111101100010000",
    "1111111111000101",
    "1111100111101001",
    "1111001001000010",
    "1110101010110010",
    "1110010011101111",
    "1110001001011101",
    "1110001110001101",
    "1110011110011001",
    "1110110010111011",
    "1111000101000101",
    "1111010000110000",
    "1111010110010010",
    "1111011000010000",
    "1111011001011000",
    "1111011100011110",
    "1111100100001110",
    "1111110001111110",
    "1111111010010001",
    "1111100010100001",
    "1111001001111101",
    "1110110011110100",
    "1110100010101001",
    "1110011000100101",
    "1110010110011000",
    "1110011010101000",
    "1110100010010101",
    "1110101010001001",
    "1110101111111111",
    "1110110011000000",
    "1110110011010101",
    "1110110010011100",
    "1110110010111011",
    "1110110111000110",
    "1111000000000011",
    "1111001101001100",
    "1111011100100101",
    "1111101100001111",
    "1111111010101100",
    "1111111000100011",
    "1111101101011111",
    "1111100011111011",
    "1111011011100110",
    "1111010100101001",
    "1111001111011111",
    "1111001100010011",
    "1111001010100011",
    "1111001001000110",
    "1111000110101101",
    "1111000011001000",
    "1110111111001010",
    "1110111100010001",
    "1110111011101011",
    "1110111101111010",
    "1111000010110100",
    "1111001001101101",
    "1111010001100010",
    "1111011001011001",
    "1111100000110110",
    "1111101001001010",
    "1111110101101100",
    "1111110110101001",
    "1111011011110000",
    "1110111100011100",
    "1110011110001001",
    "1110000110101101",
    "1101111010110100",
    "1101111100010011",
    "1110001000101101",
    "1110011010011001",
    "1110101011101101",
    "1110111000100000",
    "1110111111010111",
    "1111000001100100",
    "1111000001100001",
    "1111000001110000",
    "1111000100000011",
    "1111001000001000",
    "1111001100100000",
    "1111001111100100",
    "1111010000000011",
    "1111001101111111",
    "1111001010010100",
    "1111000110000000",
    "1111000001100110",
    "1110111101010110",
    "1110111011010110",
    "1110111111111011",
    "1111001110001100",
    "1111100110011011",
    "1111111010011001",
    "1111011010100110",
    "1111000000110011",
    "1110110010011101",
    "1110110001110110",
    "1110111100100110",
    "1111001111010001",
    "1111100111110001",
    "1111111011011101",
    "1111011011101000",
    "1110111010111000",
    "1110011101000000",
    "1110000101111001",
    "1101111001011001",
    "1101111001111100",
    "1110000110001101",
    "1110011010001011",
    "1110110001000011",
    "1111001000000001",
    "1111100000010010",
    "1111111100101111",
    "1111100000110110",
    "1110111001110010",
    "1110010011011000",
    "1101110100111100",
    "1101100100101110",
    "1101100101011010",
    "1101110100011101",
    "1110001011100001",
    "1110100011100100",
    "1110110111010000",
    "1111000100110011",
    "1111001111010111",
    "1111011101011001",
    "1111110011111011",
    "1111101100000011",
    "1111000111000011",
    "1110100101001001",
    "1110001110100100",
    "1110001001000010",
    "1110010101010010",
    "1110101101011110",
    "1111001001011001",
    "1111100010000101",
    "1111110011010000",
    "1111111100011011",
    "1111111110111010",
    "1111111100000110",
    "1111110101110110",
    "1111101101000110",
    "1111100010010101",
    "1111010110110111",
    "1111001100010001",
    "1111000100111100",
    "1111000100110011",
    "1111001111010111",
    "1111100101101110",
    "1111111010110111",
    "1111011000001001",
    "1110111000011010",
    "1110100001001101",
    "1110010110100000",
    "1110011001100010",
    "1110101000001001",
    "1110111110001100",
    "1111010110111100",
    "1111101101110010",
    "1111111111011100",
    "1111110101101110",
    "1111110001011101",
    "1111110001011011",
    "1111110010110000",
    "1111110011000011",
    "1111110001011110",
    "1111110000010010",
    "1111110011110011",
    "1111111111100100",
    "1111101011010111",
    "1111001111101011",
    "1110110010110011",
    "1110011011000100",
    "1110001101101110",
    "1110001100100110",
    "1110010101001011",
    "1110100010101011",
    "1110110001000010",
    "1110111111101001",
    "1111010001000111",
    "1111100111110001",
    "1111111100100001",
    "1111011111010110",
    "1111000110110110",
    "1110111010000001",
    "1110111101111010",
    "1111010010111001",
    "1111110100011000",
    "1111100101001110",
    "1111000010000000",
    "1110100111101101",
    "1110011001010000",
    "1110010111001101",
    "1110011111111000",
    "1110110000000010",
    "1111000011111100",
    "1111010111111100",
    "1111101000100100",
    "1111110011001000",
    "1111110101110111",
    "1111110000001000",
    "1111100011000001",
    "1111010001111011",
    "1111000001010100",
    "1110110101010011",
    "1110110000010001",
    "1110110010011010",
    "1110111010000010",
    "1111000011101001",
    "1111001011011001",
    "1111001110100001",
    "1111001100101110",
    "1111001001101111",
    "1111001010111111",
    "1111010100011010",
    "1111100111000101",
    "1111111111100000",
    "1111100100011101",
    "1111001101010100",
    "1110111110101101",
    "1110111010001011",
    "1110111101110000",
    "1111000110010000",
    "1111010000100110",
    "1111011010100011",
    "1111100100000110",
    "1111101111111111",
    "1111111110001001",
    "1111100100101001",
    "1111000101011111",
    "1110100110011011",
    "1110001110100110",
    "1110000100000011",
    "1110001001101111",
    "1110011101000100",
    "1110110111100101",
    "1111010010000011",
    "1111100110110001",
    "1111110010100011",
    "1111110101111110",
    "1111110101100100",
    "1111111000010010",
    "1111111100110100",
    "1111101001010010",
    "1111010001000010",
    "1110111010100011",
    "1110101100001111",
    "1110101010000100",
    "1110110100000001",
    "1111001000000100",
    "1111100011110110",
    "1111111011110100",
    "1111011011000001",
    "1110111110010111",
    "1110101011000010",
    "1110100110000001",
    "1110110011100111",
    "1111010100101010",
    "1111111011011001",
    "1111000101001110",
    "1110010011001011",
    "1101101110011110",
    "1101011100100110",
    "1101011110011001",
    "1101101111000000",
    "1110000110010101",
    "1110011111100011",
    "1110111010100101",
    "1111011000111111",
    "1111111011100100",
    "1111100000011100",
    "1111000000100011",
    "1110101010001111",
    "1110100001011100",
    "1110100101111001",
    "1110110010110011",
    "1111000010001111",
    "1111001111000101",
    "1111010110101101",
    "1111011010000001",
    "1111011011011001",
    "1111011101010010",
    "1111100001011100",
    "1111100111100001",
    "1111101101101000",
    "1111110011010010",
    "1111111010011111",
    "1111111001011110",
    "1111100110100101",
    "1111001101101110",
    "1110110011100010",
    "1110011110011111",
    "1110010100010010",
    "1110010111000001",
    "1110100011110100",
    "1110110100110011",
    "1111000101101110",
    "1111010101101110",
    "1111100110001001",
    "1111111000111001",
    "1111110001011011",
    "1111011010011000",
    "1111000101011000",
    "1110110110111011",
    "1110110010000010",
    "1110110110001011",
    "1111000000010111",
    "1111001101010110",
    "1111011011010001",
    "1111101010010101",
    "1111111011011101",
    "1111110000110001",
    "1111011011010110",
    "1111000111001011",
    "1110111000111100",
    "1110110101110110",
    "1111000001011010",
    "1111011011001010",
    "1111111110011001",
    "1111011100001001",
    "1110111100001010",
    "1110100111011111",
    "1110100001000111",
    "1110101000001011",
    "1110111001100101",
    "1111010010111110",
    "1111110010110011",
    "1111101000101110",
    "1111000010010111",
    "1110011110101000",
    "1110000010011101",
    "1101110001110100",
    "1101101110010010",
    "1101110101101010",
    "1110000011000101",
    "1110010001000011",
    "1110011011010011",
    "1110100010011101",
    "1110101011110111",
    "1110111100110000",
    "1111010111110101",
    "1111111010111100",
    "1111100000110110",
    "1111000011010111",
    "1110110010111000",
    "1110110001100001",
    "1110111011010100",
    "1111001001101101",
    "1111010110101101",
    "1111011111000010",
    "1111100011011010",
    "1111100111010101",
    "1111101111010100",
    "1111111110111010",
    "1111101010001100",
    "1111010000011111",
    "1110111010001111",
    "1110101101101000",
    "1110101110101011",
    "1110111101011110",
    "1111010110001001",
    "1111110011000000",
    "1111110001100110",
    "1111011100000111",
    "1111001111011110",
    "1111001101011100",
    "1111010110001101",
    "1111101000010001",
    "1111111111000001",
    "1111100011010000",
    "1111000111111001",
    "1110101111101011",
    "1110011100100101",
    "1110001111110011",
    "1110001001110100",
    "1110001010001111",
    "1110010000001100",
    "1110011010101011",
    "1110101000101000",
    "1110111001100111",
    "1111001111010001",
    "1111101011010101",
    "1111110010101110",
    "1111001110000010",
    "1110101011110011",
    "1110010001100100",
    "1110000011011000",
    "1110000011010101",
    "1110001111100100",
    "1110100011001000",
    "1110111000001000",
    "1111001001111100",
    "1111011001000010",
    "1111101001101101",
    "1111111111010010",
    "1111100101011010",
    "1111000111101100",
    "1110101101111000",
    "1110011101110101",
    "1110011100100101",
    "1110101100111111",
    "1111001100111000",
    "1111110110010110",
    "1111011110100011",
    "1110111001111101",
    "1110100001010111",
    "1110011000000100",
    "1110011110101000",
    "1110110000101110",
    "1111000111110100",
    "1111011110100110",
    "1111110010001011",
    "1111111100111101",
    "1111101100110100",
    "1111011100011100",
    "1111001011111101",
    "1110111011111111",
    "1110101110011011",
    "1110100101011010",
    "1110100010010101",
    "1110100101010101",
    "1110101100100001",
    "1110110101011111",
    "1110111110011100",
    "1111000110011010",
    "1111001101010100",
    "1111010011100110",
    "1111011001001110",
    "1111011111111000",
    "1111101011100010",
    "1111111111000010",
    "1111100101110100",
    "1111000110111001",
    "1110101011001110",
    "1110011001100010",
    "1110010110011010",
    "1110100010101110",
    "1110111001001011",
    "1111010001001100",
    "1111100011001000",
    "1111101011001101",
    "1111101100110010",
    "1111101110111000",
    "1111110111000110",
    "1111110111101110",
    "1111100000000011",
    "1111001000101010",
    "1110111000101010",
    "1110110101100010",
    "1110111111100100",
    "1111010001010100",
    "1111100101001101",
    "1111111001000010",
    "1111110010000111",
    "1111011001111010",
    "1110111110001111",
    "1110100010010101",
    "1110001011010001",
    "1110000000011001",
    "1110001000011011",
    "1110100100110001",
    "1111010000111000",
    "1111111100010111",
    "1111001110000000",
    "1110101100100011",
    "1110011100000001",
    "1110011011011110",
    "1110100101111011",
    "1110110101010000",
    "1111000100011111",
    "1111010010000110",
    "1111100001010111",
    "1111110110001100",
    "1111101110011011",
    "1111001110110110",
    "1110110000010100",
    "1110011000011110",
    "1110001011100001",
    "1110001011111000",
    "1110011000110100",
    "1110101111000111",
    "1111001010110111",
    "1111101000010000",
    "1111111011100111",
    "1111100010111000",
    "1111001111011110",
    "1111000010101100",
    "1110111101000100",
    "1110111110001111",
    "1111000101010011",
    "1111010001101110",
    "1111100100000011",
    "1111111100100101",
    "1111100101101010",
    "1111000101010111",
    "1110100110001001",
    "1110001100010111",
    "1101111011110000",
    "1101110110010011",
    "1101111011001001",
    "1110000110111111",
    "1110010101101110",
    "1110100011110001",
    "1110101111010100",
    "1110111000010000",
    "1110111111010010",
    "1111000101010010",
    "1111001011101111",
    "1111010101000110",
    "1111100011010000",
    "1111110101110111",
    "1111110101101101",
    "1111100011111011",
    "1111011001101011",
    "1111011011001001",
    "1111101010000110",
    "1111111011011100",
    "1111011011000010",
    "1110111011101011",
    "1110100100000000",
    "1110011000010001",
    "1110011010001011",
    "1110101010111100",
    "1111001010100000",
    "1111110101100010",
    "1111011001110111",
    "1110101011100011",
    "1110000111011000",
    "1101110011000001",
    "1101110001011001",
    "1110000000100111",
    "1110011001111010",
    "1110110100111110",
    "1111001010101010",
    "1111010111001110",
    "1111011010111101",
    "1111011000010101",
    "1111010100110011",
    "1111011000010000",
    "1111100111100000",
    "1111111101011011",
    "1111011011010100",
    "1110111010101010",
    "1110100011010111",
    "1110011010011001",
    "1110100000100111",
    "1110110001110110",
    "1111000111101111",
    "1111011100101011",
    "1111101100111001",
    "1111111000110101",
    "1111111011011011",
    "1111101100001001",
    "1111010111010101",
    "1110111110100011",
    "1110100110100010",
    "1110010100010000",
    "1110001011011001",
    "1110001101001110",
    "1110010111000011",
    "1110100011110100",
    "1110110000001101",
    "1110111101000101",
    "1111001101110101",
    "1111100100101110",
    "1111111110111110",
    "1111100001000000",
    "1111000110011011",
    "1110110100101100",
    "1110101111001010",
    "1110110101010000",
    "1111000010111001",
    "1111010011011100",
    "1111100100101110",
    "1111110111111111",
    "1111110000101000",
    "1111010101001000",
    "1110111000010000",
    "1110011111101001",
    "1110010001101110",
    "1110010010111110",
    "1110100011011100",
    "1110111110001101",
    "1111011011110011",
    "1111110100111001",
    "1111111010100001",
    "1111110001101111",
    "1111101101011010",
    "1111101010011101",
    "1111101000010000",
    "1111101001010100",
    "1111110001100111",
    "1111111011100111",
    "1111011110001100",
    "1110111010001111",
    "1110010111010101",
    "1101111101001111",
    "1101110000011100",
    "1101110000100110",
    "1101111010101000",
    "1110001100000010",
    "1110100100000011",
    "1111000010101011",
    "1111100111011000",
    "1111101111101111",
    "1111000110101100",
    "1110100010100111",
    "1110001000101100",
    "1101111100000111",
    "1101111101010111",
    "1110001010101010",
    "1110100000101110",
    "1110111011101111",
    "1111010111111111",
    "1111110010000001",
    "1111111001001100",
    "1111101100010101",
    "1111101001101001",
    "1111110001110101",
    "1111111100100000",
    "1111100100101111",
    "1111001011101011",
    "1110110110010010",
    "1110101000001100",
    "1110100010101001",
    "1110100100010101",
    "1110101010100110",
    "1110110010110110",
    "1110111011001100",
    "1111000010101001",
    "1111001001100000",
    "1111010001111001",
    "1111011111011110",
    "1111110101010100",
    "1111101011111011",
    "1111000111010110",
    "1110100010101111",
    "1110000100110111",
    "1101110011010010",
    "1101110000110001",
    "1101111100100001",
    "1110010010011111",
    "1110101101101001",
    "1111001001001011",
    "1111100001111011",
    "1111111000000010",
    "1111110001100111",
    "1111011000010000",
    "1110111011000100",
    "1110011100110000",
    "1110000010101110",
    "1101110010011101",
    "1101101111101110",
    "1101111010101000",
    "1110001110110110",
    "1110100110001101",
    "1110111010111101",
    "1111001001100010",
    "1111010001000011",
    "1111010010011001",
    "1111010001101001",
    "1111010110000000",
    "1111100100011101",
    "1111111101110000",
    "1111100001111000",
    "1111000001111110",
    "1110101001110100",
    "1110011110011111",
    "1110100001010111",
    "1110101110101000",
    "1110111111110101",
    "1111001110111010",
    "1111010111010011",
    "1111010111110100",
    "1111010010000101",
    "1111001000110100",
    "1111000001000111",
    "1111000001000011",
    "1111001100101000",
    "1111100100100100",
    "1111111010010011",
    "1111010110011010",
    "1110110110010010",
    "1110011111010111",
    "1110010100110111",
    "1110010110001011",
    "1110011111011110",
    "1110101011110000",
    "1110110110011000",
    "1110111101001110",
    "1111000001000011",
    "1111000101111100",
    "1111010001000010",
    "1111100100101100",
    "1111111111001001",
    "1111100100100100",
    "1111001100110111",
    "1110111110111011",
    "1110111101000000",
    "1111000100110011",
    "1111010000011111",
    "1111011010101000",
    "1111100000101110",
    "1111100011100010",
    "1111100101110001",
    "1111101001010110",
    "1111101110010111",
    "1111110011001100",
    "1111110100111101",
    "1111110001001010",
    "1111100111101000",
    "1111011010100000",
    "1111001101000000",
    "1111000010000011",
    "1110111011000001",
    "1110110111100011",
    "1110110111010101",
    "1110111011000100",
    "1111000100101010",
    "1111010110011011",
    "1111110001000011",
    "1111101101100000",
    "1111001001110100",
    "1110101001101011",
    "1110010010010000",
    "1110000110010101",
    "1110000101011111",
    "1110001100101010",
    "1110010111101000",
    "1110100010111011",
    "1110101100011100",
    "1110110011101110",
    "1110111001011001",
    "1110111110101000",
    "1111000100001101",
    "1111001010011001",
    "1111010000110011",
    "1111010110111110",
    "1111011100110101",
    "1111100011000000",
    "1111101011010010",
    "1111110111100000",
    "1111110111101100",
    "1111100011110100",
    "1111001111111011",
    "1110111111010010",
    "1110110100001101",
    "1110101111101000",
    "1110110000100011",
    "1110110100100100",
    "1110111001001110",
    "1110111100111100",
    "1110111111001010",
    "1111000000001010",
    "1111000000011001",
    "1111000000100001",
    "1111000001010100",
    "1111000011011000",
    "1111000110110110",
    "1111001011100000",
    "1111010000110001",
    "1111010110100101",
    "1111011111000100",
    "1111101100111011",
    "1111111110111001",
    "1111100110001101",
    "1111001101010110",
    "1110111001110010",
    "1110101111111011",
    "1110110010000010",
    "1110111110001100",
    "1111001111000100",
    "1111011110111111",
    "1111101001101000",
    "1111101101100001",
    "1111101100111111",
    "1111101101110000",
    "1111110101111010",
    "1111110111011011",
    "1111011100001100",
    "1110111110010111",
    "1110100101001001",
    "1110010111010011",
    "1110011010100011",
    "1110110000100111",
    "1111010101110110",
    "1111111100101010",
    "1111001111110101",
    "1110101011111101",
    "1110010110011111",
    "1110010001111000",
    "1110011011110011",
    "1110101110010111",
    "1111000101101010",
    "1111100000110000",
    "1111111111011011",
    "1111011110110001",
    "1110111101001010",
    "1110100001000010",
    "1110001111000111",
    "1110001011000001",
    "1110010110101100",
    "1110110001010000",
    "1111010111011000",
    "1111111100110111",
    "1111010011010010",
    "1110110010101001",
    "1110011111010100",
    "1110011010100011",
    "1110100001110001",
    "1110101111101110",
    "1110111110111010",
    "1111001011000110",
    "1111010010101110",
    "1111010110101111",
    "1111011001000111",
    "1111011011110111",
    "1111100001001010",
    "1111101011101110",
    "1111111101011001",
    "1111101010000100",
    "1111001101010111",
    "1110110000101001",
    "1110011000110000",
    "1110001010000110",
    "1110000111111100",
    "1110010011010111",
    "1110101001101101",
    "1111000101100111",
    "1111100000111011",
    "1111110110100010",
    "1111111100011010",
    "1111111000111000",
    "1111111110000100",
    "1111110110101010",
    "1111101011000111",
    "1111100110001000",
    "1111101100010101",
    "1111111110010101",
    "1111100111101011",
    "1111001100100011",
    "1110110111011000",
    "1110101101111111",
    "1110110001111101",
    "1110111111101110",
    "1111010010011010",
    "1111100110110001",
    "1111111011101111",
    "1111101110001111",
    "1111010111110101",
    "1111000011001101",
    "1110110010111101",
    "1110101010001011",
    "1110101011000110",
    "1110110101010000",
    "1111000101110001",
    "1111010111111010",
    "1111100110110001",
    "1111101111000101",
    "1111110000001010",
    "1111101011010110",
    "1111100010111101",
    "1111011001011001",
    "1111010000111001",
    "1111001011010110",
    "1111001001101111",
    "1111001100000101",
    "1111010001110000",
    "1111011001101111",
    "1111100011010011",
    "1111101110010001",
    "1111111010010101",
    "1111111000101100",
    "1111101011001001",
    "1111011101101101",
    "1111010001101001",
    "1111001000001110",
    "1111000010001011",
    "1110111111000111",
    "1110111101110111",
    "1110111101010110",
    "1110111100101000",
    "1110111011000111",
    "1110111000111010",
    "1110110110111011",
    "1110110111001000",
    "1110111101001110",
    "1111001101100000",
    "1111101001101000",
    "1111110000100101",
    "1111000111011010",
    "1110100011001101",
    "1110001011010001",
    "1110000011110001",
    "1110001100010100",
    "1110011111001010",
    "1110110100101111",
    "1111000110101111",
    "1111010010011100",
    "1111011011011000",
    "1111100111101000",
    "1111111011011010",
    "1111101000011010",
    "1111001000000011",
    "1110101010101101",
    "1110010110111001",
    "1110010000111101",
    "1110011001110010",
    "1110101111010111",
    "1111001101111010",
    "1111110000110000",
    "1111101100110000",
    "1111001111000111",
    "1110111010010011",
    "1110110000111011",
    "1110110011001000",
    "1110111110011100",
    "1111001110110101",
    "1111100010000010",
    "1111111000001011",
    "1111101110010111",
    "1111010010111000",
    "1110111000011011",
    "1110100011001000",
    "1110011000110100",
    "1110100000011001",
    "1110111101000111",
    "1111101011101100",
    "1111011100110000",
    "1110101000000100",
    "1110000000101011",
    "1101101100100001",
    "1101101011111101",
    "1101111001100000",
    "1110001101000010",
    "1110011111111010",
    "1110101110100110",
    "1110111011010110",
    "1111001100011011",
    "1111100110101000",
    "1111110101000101",
    "1111001011000010",
    "1110100011001010",
    "1110000100110001",
    "1101110101001000",
    "1101110101000101",
    "1101111111101001",
    "1110001101100110",
    "1110011001010101",
    "1110100000101001",
    "1110100101000101",
    "1110101001010000",
    "1110101110110011",
    "1110110110100000",
    "1110111111101110",
    "1111001000100010",
    "1111001111010001",
    "1111010100001000",
    "1111011010011011",
    "1111100110011010",
    "1111111010010100",
    "1111101011010101",
    "1111001111101001",
    "1110111000100101",
    "1110101010110101",
    "1110101000100000",
    "1110101111101100",
    "1110111100000101",
    "1111001001101010",
    "1111010101101010",
    "1111011111000111",
    "1111100101100000",
    "1111101000010010",
    "1111100111000111",
    "1111100001111001",
    "1111011001001011",
    "1111001111000111",
    "1111000110100111",
    "1111000010000110",
    "1111000011000101",
    "1111001001110101",
    "1111010101001101",
    "1111100011101110",
    "1111110101011000",
    "1111110100110000",
    "1111011010000001",
    "1110111011101111",
    "1110011110010110",
    "1110000111100010",
    "1101111100001111",
    "1101111110101000",
    "1110001100001100",
    "1110011111000111",
    "1110110000111101",
    "1110111100101000",
    "1111000001010000",
    "1111000011111100",
    "1111001100010110",
    "1111100000010001",
    "1111111111011000",
    "1111010111111001",
    "1110110001111001",
    "1110010110000001",
    "1110001010010011",
    "1110001110101001",
    "1110011101001110",
    "1110101110011110",
    "1110111100100110",
    "1111000111011000",
    "1111010011101110",
    "1111100110100110",
    "1111111101101000",
    "1111011011000010",
    "1110111000001110",
    "1110011100101110",
    "1110001110100011",
    "1110001111111111",
    "1110011101011001",
    "1110101111111111",
    "1111000001011111",
    "1111001111001000",
    "1111011010101011",
    "1111100111101000",
    "1111111000001010",
    "1111110011100110",
    "1111011110100011",
    "1111001101110101",
    "1111000110100000",
    "1111001011101000",
    "1111011101000101",
    "1111110111100100",
    "1111101010000110",
    "1111001101001111",
    "1110110101110111",
    "1110100110110010",
    "1110100010000011",
    "1110101001000100",
    "1110111100000100",
    "1111011001110000",
    "1111111111010111",
    "1111010111101000",
    "1110110000101001",
    "1110010000100111",
    "1101111011010001",
    "1101110010000010",
    "1101110100000000",
    "1101111110101110",
    "1110001111101001",
    "1110100110101111",
    "1111000101100100",
    "1111101100001001",
    "1111100111101000",
    "1110111010111010",
    "1110010100100010",
    "1101111010011110",
    "1101110000010100",
    "1101110101000001",
    "1110000011001111",
    "1110010100110001",
    "1110100100101010",
    "1110110010110100",
    "1111000100000000",
    "1111011100010110",
    "1111111100110110",
    "1111011101100001",
    "1110111010000110",
    "1110100000010001",
    "1110010101000001",
    "1110011010000100",
    "1110101101110101",
    "1111001100110101",
    "1111110010011100",
    "1111100110010011",
    "1111000010010100",
    "1110100110010101",
    "1110010110011111",
    "1110010100110001",
    "1110011111111011",
    "1110110011011111",
    "1111001010011001",
    "1111100001100100",
    "1111111000010100",
    "1111110001001000",
    "1111011011101010",
    "1111001000101100",
    "1110111001101011",
    "1110110000011001",
    "1110101110000111",
    "1110110001110100",
    "1110111000101100",
    "1110111111100001",
    "1111000100001010",
    "1111000110010011",
    "1111000111101100",
    "1111001010100101",
    "1111001111111011",
    "1111011000011011",
    "1111100101001110",
    "1111110111000001",
    "1111110011001101",
    "1111011100010110",
    "1111001000011110",
    "1110111011110000",
    "1110111001010101",
    "1111000010011101",
    "1111010100110110",
    "1111101010111000",
    "1111111110011011",
    "1111110101011100",
    "1111110010110101",
    "1111111001001100",
    "1111111010001001",
    "1111101101011101",
    "1111100111111111",
    "1111101110001011",
    "1111111111100110",
    "1111100101110100",
    "1111001011100110",
    "1110110111101000",
    "1110101110011001",
    "1110110000100110",
    "1110111011001110",
    "1111001001110101",
    "1111011001001001",
    "1111101000111000",
    "1111111010111100",
    "1111101111101000",
    "1111011000011110",
    "1111000011110011",
    "1110110111000100",
    "1110110110011111",
    "1111000010100111",
    "1111010111110001",
    "1111101111001101",
    "1111111101110011",
    "1111110011110110",
    "1111110011101010",
    "1111111010101001",
    "1111111011001001",
    "1111110001010101",
    "1111101010010001",
    "1111100111010111",
    "1111101001010110",
    "1111110000001000",
    "1111111010101001",
    "1111111000101101",
    "1111101011101001",
    "1111011111110110",
    "1111010111001011",
    "1111010011001111",
    "1111010100100101",
    "1111011010111100",
    "1111100101010101",
    "1111110010010011",
    "1111111111110000",
    "1111110100111010",
    "1111101110001011",
    "1111101101101000",
    "1111110011011001",
    "1111111101110010",
    "1111110110001110",
    "1111101100101101",
    "1111101001001111",
    "1111101101110011",
    "1111111010001000",
    "1111110100011110",
    "1111100010101110",
    "1111010110000000",
    "1111010011001010",
    "1111011100111111",
    "1111110011001000",
    "1111101101110111",
    "1111001011101111",
    "1110101100101011",
    "1110010101110001",
    "1110001001111001",
    "1110001001001001",
    "1110010001011001",
    "1110011111001111",
    "1110101111000000",
    "1110111110111111",
    "1111010000111001",
    "1111100111011010",
    "1111111100011110",
    "1111011100110011",
    "1110111110101011",
    "1110100111111001",
    "1110011100111010",
    "1110011111010110",
    "1110101011111111",
    "1110111100010100",
    "1111001010001100",
    "1111010001100001",
    "1111010011000101",
    "1111010101100000",
    "1111100000011010",
    "1111111000000000",
    "1111100101001000",
    "1110111110111000",
    "1110011111011001",
    "1110001111000000",
    "1110010001111101",
    "1110100101001011",
    "1111000000001100",
    "1111011010001011",
    "1111101100110111",
    "1111110110011000",
    "1111111000010111",
    "1111110101010001",
    "1111101111110011",
    "1111101010000010",
    "1111100100000101",
    "1111011101101110",
    "1111011000011000",
    "1111010111000011",
    "1111011101001111",
    "1111101100100110",
    "1111111100011110",
    "1111100010101011",
    "1111001011111010",
    "1110111101001100",
    "1110111000111100",
    "1110111110111000",
    "1111001101100000",
    "1111100010100110",
    "1111111011111010",
    "1111101001001001",
    "1111010000011100",
    "1110111110001001",
    "1110110101100010",
    "1110111000001011",
    "1111000100010011",
    "1111010110000110",
    "1111101010110111",
    "1111111110100010",
    "1111100110111010",
    "1111001111000101",
    "1110111001000111",
    "1110100111100011",
    "1110011100111010",
    "1110011011110111",
    "1110100100110111",
    "1110110100110111",
    "1111000110111110",
    "1111010101110110",
    "1111011101111111",
    "1111011111000100",
    "1111011011000010",
    "1111010101001011",
    "1111010000101011",
    "1111001110101000",
    "1111001110011001",
    "1111001110011111",
    "1111001101010010",
    "1111001001101101",
    "1111000011100001",
    "1110111011001110",
    "1110110001100001",
    "1110100111011010",
    "1110011110100011",
    "1110011001101111",
    "1110011100100101",
    "1110101001110000",
    "1111000001101110",
    "1111100010010000",
    "1111111001000100",
    "1111010101100010",
    "1110110111111001",
    "1110100011010011",
    "1110011000011010",
    "1110010101110010",
    "1110011001000111",
    "1110100000010100",
    "1110101001111100",
    "1110110100111011",
    "1111000000000011",
    "1111001010000100",
    "1111010001011111",
    "1111010101001000",
    "1111010100101111",
    "1111010001011100",
    "1111001101001111",
    "1111001010000111",
    "1111001001000110",
    "1111001010000111",
    "1111001100000100",
    "1111001101100110",
    "1111001110101001",
    "1111010001001010",
    "1111010111111010",
    "1111100100101010",
    "1111110111000001",
    "1111110011111000",
    "1111100000000000",
    "1111010000110000",
    "1111000111100011",
    "1111000011010011",
    "1111000001000011",
    "1110111101111010",
    "1110111000101100",
    "1110110010110110",
    "1110101111010110",
    "1110110001001111",
    "1110111010010001",
    "1111001001111001",
    "1111011101100001",
    "1111110010000000",
    "1111111010111100",
    "1111101010000110",
    "1111011010111010",
    "1111001100111101",
    "1111000000100001",
    "1110110110110100",
    "1110110001100001",
    "1110110001101011",
    "1110110111000001",
    "1111000000100001",
    "1111001110000101",
    "1111100000011111",
    "1111110111110100",
    "1111101101011010",
    "1111010010100110",
    "1110111011111111",
    "1110101101011100",
    "1110101001001001",
    "1110101110010110",
    "1110111001000100",
    "1111000101001101",
    "1111010010000000",
    "1111100001010111",
    "1111110101011100",
    "1111110001010010",
    "1111010101100101",
    "1110111100010100",
    "1110101011000001",
    "1110100110001110",
    "1110101110000111",
    "1110111110001101",
    "1111010000001000",
    "1111011101101000",
    "1111100011010011",
    "1111100001101100",
    "1111011011011110",
    "1111010100010000",
    "1111001110110101",
    "1111001100100000",
    "1111001111000111",
    "1111011000101000",
    "1111101001011011",
    "1111111111110010",
    "1111100110010110",
    "1111001110101110",
    "1110111101100100",
    "1110110110010110",
    "1110111001001001",
    "1111000010001010",
    "1111001011111100",
    "1111010011001000",
    "1111011000111010",
    "1111100001001000",
    "1111101110111010",
    "1111111101011100",
    "1111100111010101",
    "1111010100100111",
    "1111001011011000",
    "1111001111001100",
    "1111011110010111",
    "1111110010100100",
    "1111111011101011",
    "1111110001110011",
    "1111101110101010",
    "1111101100000000",
    "1111100011111011",
    "1111010011110011",
    "1110111110001010",
    "1110101001110000",
    "1110011101111000",
    "1110011111110110",
    "1110110000110110",
    "1111001101010100",
    "1111101111011101",
    "1111101110010110",
    "1111001111110001",
    "1110110110010011",
    "1110100011000001",
    "1110010110111011",
    "1110010010011100",
    "1110010101111100",
    "1110100001111101",
    "1110110110011000",
    "1111010001110011",
    "1111110001001110",
    "1111101111011000",
    "1111010011110011",
    "1110111110001101",
    "1110101111010010",
    "1110100110110001",
    "1110100011101110",
    "1110100100111001",
    "1110101000110111",
    "1110101110011100",
    "1110110100101010",
    "1110111010101010",
    "1110111111110000",
    "1111000011110001",
    "1111000110101111",
    "1111001001000100",
    "1111001011000111",
    "1111001100111000",
    "1111001110001100",
    "1111001110011111",
    "1111001101010010",
    "1111001001111111",
    "1111000100100000",
    "1110111101100100",
    "1110110110111111",
    "1110110100101010",
    "1110111011010100",
    "1111001101110010",
    "1111101011101101",
    "1111101110100101",
    "1111000111011111",
    "1110100101110001",
    "1110001111001101",
    "1110000110011011",
    "1110001001101010",
    "1110010100100100",
    "1110100010100100",
    "1110110000000010",
    "1110111011010110",
    "1111000100001011",
    "1111001010101010",
    "1111010000001000",
    "1111011000001011",
    "1111100110011111",
    "1111111100100011",
    "1111100111010001",
    "1111001010000001",
    "1110110001101100",
    "1110100011011000",
    "1110100010100010",
    "1110101110001010",
    "1111000000111000",
    "1111010100000110",
    "1111100001110001",
    "1111101000101101",
    "1111101101100111",
    "1111110110000010",
    "1111111010000000",
    "1111100010011100",
    "1111001000010110",
    "1110110011100110",
    "1110101101000010",
    "1110111010100101",
    "1111011010011000",
    "1111111011111100",
    "1111010011111000",
    "1110110111101101",
    "1110101100111111",
    "1110110011111011",
    "1111001001000111",
    "1111100111110010",
    "1111110100010001",
    "1111001110100001",
    "1110101001111101",
    "1110001010000010",
    "1101110010001111",
    "1101100101101010",
    "1101100101111110",
    "1101110001001100",
    "1110000010000000",
    "1110010010101110",
    "1110011111011001",
    "1110101000010110",
    "1110110010011001",
    "1111000011000001",
    "1111011101110010",
    "1111111110000011",
    "1111010110100101",
    "1110110011111001",
    "1110011101000010",
    "1110010101110001",
    "1110011100011011",
    "1110101011101010",
    "1110111101101000",
    "1111001110001100",
    "1111011011110000",
    "1111100110100010",
    "1111101111000101",
    "1111110101110010",
    "1111111100000101",
    "1111111011001010",
    "1111101101011010",
    "1111011001011000",
    "1111000000110001",
    "1110101000011010",
    "1110010101110001",
    "1110001101111101",
    "1110010011101100",
    "1110100100110011",
    "1110111100101101",
    "1111010111110010",
    "1111110011110000",
    "1111110000011010",
    "1111010101110001",
    "1110111110011100",
    "1110101101001010",
    "1110100101101111",
    "1110101100000010",
    "1111000000100111",
    "1111100000000000",
    "1111111011110100",
    "1111011010000100",
    "1111000000110110",
    "1110110011111000",
    "1110110100101010",
    "1111000010101111",
    "1111011011111100",
    "1111111100111001",
    "1111011111000000",
    "1110111101001010",
    "1110100010011010",
    "1110010010011111",
    "1110001111001000",
    "1110010111010001",
    "1110100111010001",
    "1110111010011001",
    "1111001100011100",
    "1111011010111111",
    "1111100101011101",
    "1111101100100000",
    "1111110001110000",
    "1111111000111011",
    "1111111001101001",
    "1111100011111110",
    "1111000111001011",
    "1110100111110001",
    "1110001011111000",
    "1101111000110100",
    "1101110010010111",
    "1101111001101000",
    "1110001100011110",
    "1110101000000001",
    "1111001001001100",
    "1111101100110110",
    "1111110000010101",
    "1111010010101100",
    "1110111101111111",
    "1110110100000001",
    "1110110100101100",
    "1110111101000101",
    "1111001000010110",
    "1111010001110110",
    "1111010110110010",
    "1111010110011010",
    "1111010001110110",
    "1111001011101111",
    "1111000111001011",
    "1111000110101100",
    "1111001011010001",
    "1111010100101111",
    "1111100010000010",
    "1111110000111000",
    "1111111110001101",
    "1111111000111010",
    "1111110110110111",
    "1111111100011000",
    "1111110111101000",
    "1111101000011000",
    "1111011010010100",
    "1111010010001101",
    "1111010011011100",
    "1111011111010110",
    "1111110100110000",
    "1111101111101110",
    "1111010010011100",
    "1110110111100000",
    "1110100010011001",
    "1110010101010011",
    "1110010000111110",
    "1110010100110110",
    "1110011111001101",
    "1110101110010001",
    "1110111111101110",
    "1111010010100110",
    "1111101000001011",
    "1111111110010011",
    "1111100001100111",
    "1111000100011101",
    "1110101011011000",
    "1110011010110000",
    "1110010101011011",
    "1110011011100001",
    "1110101010011001",
    "1111000000010010",
    "1111011100001100",
    "1111111100011000",
    "1111100001001111",
    "1111000000010001",
    "1110100100100000",
    "1110010000110011",
    "1110000110110110",
    "1110000101100111",
    "1110001001011001",
    "1110001110100110",
    "1110010010100100",
    "1110010100011101",
    "1110010101010011",
    "1110010110110001",
    "1110011010111100",
    "1110100100000101",
    "1110110011001011",
    "1111000111101000",
    "1111011111011010",
    "1111110111000110",
    "1111110100100011",
    "1111100101100101",
    "1111011100011110",
    "1111011000011000",
    "1111010110111111",
    "1111010101101100",
    "1111010010101011",
    "1111001101101000",
    "1111000111110111",
    "1111000010111001",
    "1110111111101110",
    "1110111111001000",
    "1111000001011001",
    "1111000101110110",
    "1111001010110000",
    "1111001101001010",
    "1111001010011110",
    "1111000010001000",
    "1110110101101110",
    "1110101000110000",
    "1110011111100110",
    "1110011101011110",
    "1110100011011101",
    "1110101111110110",
    "1110111110110011",
    "1111001101010100",
    "1111011011100000",
    "1111101100000000",
    "1111111110100010",
    "1111100011101100",
    "1111000110000000",
    "1110101010001111",
    "1110010101110010",
    "1110001100101101",
    "1110001111111011",
    "1110011100110010",
    "1110101110101000",
    "1111000000110110",
    "1111010000101110",
    "1111011101101000",
    "1111100111101010",
    "1111101111001101",
    "1111110100110100",
    "1111111001100101",
    "1111111111110010",
    "1111110110001100",
    "1111100111110100",
    "1111010110100000",
    "1111000110000011",
    "1110111011000111",
    "1110111010001011",
    "1111000101101001",
    "1111011100011011",
    "1111111010000001",
    "1111100111010001",
    "1111001100100001",
    "1110111000100111",
    "1110101100010100",
    "1110100110111001",
    "1110100110100000",
    "1110101001010000",
    "1110101101110111",
    "1110110011110011",
    "1110111010101101",
    "1111000010000010",
    "1111001000101000",
    "1111001101010100",
    "1111001111011100",
    "1111001111011100",
    "1111001110110001",
    "1111001111111011",
    "1111010101101010",
    "1111100001110011",
    "1111110100001110",
    "1111110101101000",
    "1111011111101001",
    "1111001101000100",
    "1110111111101011",
    "1110110111010000",
    "1110110010000011",
    "1110101101111010",
    "1110101000111100",
    "1110100010011111",
    "1110011011000111",
    "1110010011111011",
    "1110001101110011",
    "1110001001010000",
    "1110000110010011",
    "1110000101011011",
    "1110000111001101",
    "1110001100000101",
    "1110010100000101",
    "1110011110101001",
    "1110101011110000",
    "1110111100101101",
    "1111010010101110",
    "1111101101101011",
    "1111110100011011",
    "1111010111100010",
    "1111000000000000",
    "1110110001011001",
    "1110101101011110",
    "1110110010101110",
    "1110111100111000",
    "1111000111000100",
    "1111001110001101",
    "1111010100001010",
    "1111011101111010",
    "1111101111110011",
    "1111110100101100",
    "1111010010011100",
    "1110110000010101",
    "1110010111100000",
    "1110010000010101",
    "1110011110001010",
    "1110111101010110",
    "1111100101001011",
    "1111110100101100",
    "1111011000111010",
    "1111001011011000",
    "1111001011011101",
    "1111010110100100",
    "1111101010100100",
    "1111111010000101",
    "1111011001001100",
    "1110110101100111",
    "1110010100000000",
    "1101111001101101",
    "1101101011100110",
    "1101101100010011",
    "1101111001100010",
    "1110001101101101",
    "1110100010111110",
    "1110110100110001",
    "1111000001011110",
    "1111001001110010",
    "1111001111100110",
    "1111010101011000",
    "1111011100100101",
    "1111100100101111",
    "1111101100101111",
    "1111110100101000",
    "1111111110010101",
    "1111110011101100",
    "1111100000110011",
    "1111001011001111",
    "1110111000000011",
    "1110101100110101",
    "1110101101010100",
    "1110111001101010",
    "1111001101100110",
    "1111100010100001",
    "1111110010000100",
    "1111111000100100",
    "1111110101111110",
    "1111101110000100",
    "1111100111101011",
    "1111101001001001",
    "1111110100101110",
    "1111110111110110",
    "1111100010011001",
    "1111010001001111",
    "1111001000111111",
    "1111001010111100",
    "1111010100000001",
    "1111011111010010",
    "1111101000111011",
    "1111101110111110",
    "1111110001010111",
    "1111110001000000",
    "1111101111111000",
    "1111110010001101",
    "1111111011110100",
    "1111110010011101",
    "1111011010110000",
    "1111000001100001",
    "1110101011111000",
    "1110011110000010",
    "1110011010100000",
    "1110100001011010",
    "1110110000111110",
    "1111000110100100",
    "1111011110101011",
    "1111110101111000",
    "1111110110001001",
    "1111100110101110",
    "1111011011100001",
    "1111010011001101",
    "1111001100011110",
    "1111000110101000",
    "1111000001111011",
    "1110111111011001",
    "1111000000001000",
    "1111000100101001",
    "1111001100101110",
    "1111010111111010",
    "1111100101010101",
    "1111110011011011",
    "1111111111110000",
    "1111110110001010",
    "1111110000101111",
    "1111110000000100",
    "1111110100010100",
    "1111111100111110",
    "1111110111001110",
    "1111101010101010",
    "1111100000000010",
    "1111011001110010",
    "1111011001011101",
    "1111011111100100",
    "1111101011101111",
    "1111111100111101",
    "1111101101111101",
    "1111010110100100",
    "1110111110101000",
    "1110101000010101",
    "1110010101111100",
    "1110001001011011",
    "1110000011110011",
    "1110000100110110",
    "1110001011001111",
    "1110010101011011",
    "1110100010011100",
    "1110110010011100",
    "1111000101110111",
    "1111011100011001",
    "1111110100011001",
    "1111110100110010",
    "1111100010011010",
    "1111010111001000",
    "1111010100000000",
    "1111011000001001",
    "1111100001011100",
    "1111101101010110",
    "1111111001011001",
    "1111111100011011",
    "1111110110001011",
    "1111110101010010",
    "1111111010000000",
    "1111111100111000",
    "1111110001110011",
    "1111100111100010",
    "1111100000010111",
    "1111011101010110",
    "1111011110001101",
    "1111100001011100",
    "1111100101001000",
    "1111100111010111",
    "1111101000111000",
    "1111101110010101",
    "1111111100100000",
    "1111101010100001",
    "1111001000110111",
    "1110100100110110",
    "1110000110001110",
    "1101110011110001",
    "1101110001000000",
    "1101111011101111",
    "1110001101111000",
    "1110100000111101",
    "1110101111110101",
    "1110111000110101",
    "1110111101000100",
    "1110111110101000",
    "1111000000000010",
    "1111000011010010",
    "1111001010101010",
    "1111011000110010",
    "1111101110001010",
    "1111110111001110",
    "1111011011011011",
    "1111000011100111",
    "1110110100100000",
    "1110110001101001",
    "1110111010111101",
    "1111001100000111",
    "1111011110101000",
    "1111101100110111",
    "1111110110000101",
    "1111111110100110",
    "1111110100110010",
    "1111100001101001",
    "1111001001010001",
    "1110110001000010",
    "1110011111011100",
    "1110011001101111",
    "1110100001010100",
    "1110110010000101",
    "1111000101010011",
    "1111010111001000",
    "1111101000001000",
    "1111111011011000",
    "1111101101000100",
    "1111010010011100",
    "1110111000101101",
    "1110100101011101",
    "1110011110000101",
    "1110100100011100",
    "1110110101000011",
    "1111001001100011",
    "1111011011000100",
    "1111100100111001",
    "1111100111110010",
    "1111101001011110",
    "1111110000100101",
    "1111111110110001",
    "1111100101011011",
    "1111001000100010",
    "1110101111001000",
    "1110011111110101",
    "1110011101101101",
    "1110100110111001",
    "1110110110001101",
    "1111000110101101",
    "1111010110001110",
    "1111100100111001",
    "1111110011011000",
    "1111111110100000",
    "1111110010000101",
    "1111101001101000",
    "1111101000001000",
    "1111101111100011",
    "1111111111100000",
    "1111101011000000",
    "1111010100110001",
    "1111000010100010",
    "1110110111010110",
    "1110110100011111",
    "1110111010000010",
    "1111000111001001",
    "1111011010011101",
    "1111110010000110",
    "1111110100000010",
    "1111011010010110",
    "1111000011010000",
    "1110110000111000",
    "1110100100101110",
    "1110011111010001",
    "1110100000010010",
    "1110100111001001",
    "1110110011001101",
    "1111000011110100",
    "1111011000001000",
    "1111101110101111",
    "1111111010010101",
    "1111100101011101",
    "1111010100110100",
    "1111001010010011",
    "1111000110101100",
    "1111001001000010",
    "1111001111000010",
    "1111010110100000",
    "1111011111111111",
    "1111101110001111",
    "1111111100101000",
    "1111100001000010",
    "1111000010011010",
    "1110100110101111",
    "1110010100001011",
    "1110001111010111",
    "1110011001000010",
    "1110101101001100",
    "1111000101101001",
    "1111011101010010",
    "1111110010000110",
    "1111111011010000",
    "1111101001110001",
    "1111011001011000",
    "1111001011000100",
    "1111000001010010",
    "1110111111010010",
    "1111001000000001",
    "1111011100110000",
    "1111111011110010",
    "1111011111001100",
    "1110111010010001",
    "1110011011011001",
    "1110000111001110",
    "1110000000000111",
    "1110000101011010",
    "1110010011100100",
    "1110100101100111",
    "1110110110110001",
    "1111000100010000",
    "1111001111111000",
    "1111011110011110",
    "1111110100001101",
    "1111101101111111",
    "1111001100001110",
    "1110101110100011",
    "1110011110000010",
    "1110100001011111",
    "1110111010000110",
    "1111100001111001",
    "1111110000110011",
    "1111000111111110",
    "1110101010101011",
    "1110011011101000",
    "1110011001111100",
    "1110100010100111",
    "1110110001010010",
    "1111000010001111",
    "1111010010111011",
    "1111100001011001",
    "1111101100011010",
    "1111110011010010",
    "1111110101100101",
    "1111110011101110",
    "1111101111011000",
    "1111101011100110",
    "1111101011110010",
    "1111110010011001",
    "1111111111110100",
    "1111101100001101",
    "1111010110001110",
    "1111000010011010",
    "1110110100101010",
    "1110101111001101",
    "1110110001111110",
    "1110111010110100",
    "1111000111000100",
    "1111010101011011",
    "1111100101110001",
    "1111110111111010",
    "1111110101010010",
    "1111100100110111",
    "1111011010110000",
    "1111011010101101",
    "1111100110011000",
    "1111111011110111",
    "1111101001110010",
    "1111010000100011",
    "1110111101010100",
    "1110110010101011",
    "1110110000010010",
    "1110110011111001",
    "1110111010000111",
    "1110111111101100",
    "1111000010101110",
    "1111000010100111",
    "1110111111111101",
    "1110111011111111",
    "1110110111111001",
    "1110110100111011",
    "1110110101100101",
    "1110111101010110",
    "1111001110101001",
    "1111101000111100",
    "1111110111110110",
    "1111011010100011",
    "1111000101111110",
    "1110111111001010",
    "1111000111011101",
    "1111011011110000",
    "1111110110010010",
    "1111101111000110",
    "1111011001010011",
    "1111001010101010",
    "1111000011101001",
    "1111000011101001",
    "1111001001101101",
    "1111010101010010",
    "1111100110010011",
    "1111111100101010",
    "1111101000110100",
    "1111001100111100",
    "1110110011101010",
    "1110100000110001",
    "1110010110000100",
    "1110010010111110",
    "1110010101011011",
    "1110011100010011",
    "1110100111110111",
    "1110111000111001",
    "1111001111011100",
    "1111101010001101",
    "1111111001011110",
    "1111011111000000",
    "1111001001110000",
    "1110111011110010",
    "1110110100111100",
    "1110110011011100",
    "1110110101001101",
    "1110111000110010",
    "1110111101101011",
    "1111000100100100",
    "1111010000001111",
    "1111100100001011",
    "1111111110101111",
    "1111011011110011",
    "1110111001110010",
    "1110100000101001",
    "1110010110011010",
    "1110011101101110",
    "1110110100111100",
    "1111010110010101",
    "1111111010101110",
    "1111100100011010",
    "1111001011110011",
    "1110111101010111",
    "1110111001000110",
    "1110111101100011",
    "1111001000100111",
    "1111011000000011",
    "1111101010000001",
    "1111111110101011",
    "1111101000011101",
    "1111001011000001",
    "1110101010100101",
    "1110001011001100",
    "1101110001111011",
    "1101100010111001",
    "1101100000101011",
    "1101101010110111",
    "1101111101110011",
    "1110010110001011",
    "1110110011000000",
    "1111010100010010",
    "1111111010000010",
    "1111011101100000",
    "1110110110110010",
    "1110010110110010",
    "1110000010011111",
    "1101111100110010",
    "1110000011110100",
    "1110010100100000",
    "1110101101011100",
    "1111001101001110",
    "1111110010010111",
    "1111100101101010",
    "1110111111100100",
    "1110100000000111",
    "1110001011111100",
    "1110000110001011",
    "1110001101001111",
    "1110011100000111",
    "1110101101001001",
    "1110111011001001",
    "1111000011101010",
    "1111000110111111",
    "1111000110101010",
    "1111000100111011",
    "1111000011010000",
    "1111000001010010",
    "1110111110010110",
    "1110111010000100",
    "1110110101110001",
    "1110110101101111",
    "1110111110101101",
    "1111010010011101",
    "1111101111001000",
    "1111110000110110",
    "1111010100010111",
    "1111000000110101",
    "1110111001010000",
    "1110111100000101",
    "1111000100001010",
    "1111001011101000",
    "1111001110000010",
    "1111001001111001",
    "1111000000111011",
    "1110110101111001",
    "1110101011101011",
    "1110100100101111",
    "1110100001110100",
    "1110100010110011",
    "1110100111000110",
    "1110101110010001",
    "1110111000111110",
    "1111001001000110",
    "1111100000000011",
    "1111111101001111",
    "1111100010010111",
    "1111000011011100",
    "1110101010011011",
    "1110011010100010",
    "1110010100111110",
    "1110011000001001",
    "1110100000001111",
    "1110101000110100",
    "1110101110010111",
    "1110101111111111",
    "1110101110101101",
    "1110101100101000",
    "1110101011110111",
    "1110101101111101",
    "1110110011010101",
    "1110111011010110",
    "1111000101011011",
    "1111010010100010",
    "1111100100010011",
    "1111111011001100",
    "1111101010100011",
    "1111010001011001",
    "1110111110011100",
    "1110110101100010",
    "1110110111101111",
    "1111000010110001",
    "1111010001011111",
    "1111011101111010",
    "1111100010111011",
    "1111011110001010",
    "1111010000110001",
    "1110111110101001",
    "1110101100110010",
    "1110011111011111",
    "1110011001001011",
    "1110011010000001",
    "1110100000010100",
    "1110101001000001",
    "1110110001010101",
    "1110110111111001",
    "1110111110010100",
    "1111001000010110",
    "1111011000111110",
    "1111110000111000",
    "1111110001111101",
    "1111010100011000",
    "1110111011110101",
    "1110101100111010",
    "1110101001010000",
    "1110101110100011",
    "1110111000010110",
    "1111000010011111",
    "1111001010101010",
    "1111010000110011",
    "1111010110110111",
    "1111100000011111",
    "1111110001001100",
    "1111110110000110",
    "1111011000011000",
    "1110111011110000",
    "1110100111011010",
    "1110100001001100",
    "1110101011100011",
    "1111000100011000",
    "1111100110001000",
    "1111110101110010",
    "1111010101010000",
    "1110111100000101",
    "1110101011110111",
    "1110100100001011",
    "1110100011011111",
    "1110100111100101",
    "1110101110100001",
    "1110110110100101",
    "1110111110101001",
    "1111001000100000",
    "1111010111110100",
    "1111101110101000",
    "1111110011111100",
    "1111010100000110",
    "1110110111101111",
    "1110100100001011",
    "1110011100111100",
    "1110100001100110",
    "1110101101000111",
    "1110111001001100",
    "1111000000111001",
    "1111000011001010",
    "1111000100111100",
    "1111001101001111",
    "1111100000000101",
    "1111111100111101",
    "1111100010100110",
    "1111001000010001",
    "1110111100000111",
    "1111000010101001",
    "1111011001110111",
    "1111111001100101",
    "1111101000001011",
    "1111010011101001",
    "1111001100100001",
    "1111010001100110",
    "1111011111001010",
    "1111110000100001",
    "1111111110110110",
    "1111110001001001",
    "1111100110011110",
    "1111011101111111",
    "1111010111001110",
    "1111010100010010",
    "1111011000111010",
    "1111100111000110",
    "1111111101101010",
    "1111100111111110",
    "1111010000001111",
    "1111000001010010",
    "1110111111110001",
    "1111001100110010",
    "1111100100101111",
    "1111111110011010",
    "1111100011010111",
    "1111001111100001",
    "1111000101110110",
    "1111000110101111",
    "1111010000001100",
    "1111011110010010",
    "1111101101001001",
    "1111111001101001",
    "1111111101111110",
    "1111111001111101",
    "1111111001100010",
    "1111111010011011",
    "1111111000000110",
    "1111101101111100",
    "1111011001111010",
    "1110111101101110",
    "1110011111000000",
    "1110000100100101",
    "1101110100000101",
    "1101110000101011",
    "1101111001101010",
    "1110001011000010",
    "1110011111110110",
    "1110110011100111",
    "1111000011110110",
    "1111010000111011",
    "1111011100110111",
    "1111101001101011",
    "1111110111110101",
    "1111111010011111",
    "1111110000011001",
    "1111101100100001",
    "1111110000010100",
    "1111111010110100",
    "1111110111000101",
    "1111101000111011",
    "1111011100111010",
    "1111010011011010",
    "1111001011100101",
    "1111000100100000",
    "1110111101100001",
    "1110110110011011",
    "1110101111111000",
    "1110101010110101",
    "1110101000001000",
    "1110101000001100",
    "1110101010101101",
    "1110101110100100",
    "1110110010101111",
    "1110110110100010",
    "1110111001100111",
    "1110111011110000",
    "1110111100110010",
    "1110111100010111",
    "1110111010011000",
    "1110110110111001",
    "1110110010100010",
    "1110101110010111",
    "1110101011111100",
    "1110101101101001",
    "1110110110001110",
    "1111000111011010",
    "1111100000101100",
    "1111111110101101",
    "1111100011111001",
    "1111001100101110",
    "1110111111110000",
    "1110111101100100",
    "1111000011001010",
    "1111001011001111",
    "1111010000101100",
    "1111010000001010",
    "1111001001001100",
    "1110111101111000",
    "1110110001101001",
    "1110100111111010",
    "1110100010100100",
    "1110100001100110",
    "1110100011100111",
    "1110100110110010",
    "1110101001101000",
    "1110101011101010",
    "1110101101010001",
    "1110101111000101",
    "1110110001010010",
    "1110110011101100",
    "1110110110001110",
    "1110111000111001",
    "1110111011101000",
    "1110111110101001",
    "1111000100001011",
    "1111001111100110",
    "1111100010110011",
    "1111111100101011",
    "1111100111000001",
    "1111001110101001",
    "1110111111101100",
    "1110111101100110",
    "1111000111111111",
    "1111011010011000",
    "1111101110101111",
    "1111111111110001",
    "1111110101100001",
    "1111110001001110",
    "1111110001101001",
    "1111110100100000",
    "1111110111001100",
    "1111110111001011",
    "1111110010000000",
    "1111100110000011",
    "1111010011110011",
    "1110111101110011",
    "1110100111111001",
    "1110010110010101",
    "1110001101000111",
    "1110001110100100",
    "1110011010000110",
    "1110101011111101",
    "1110111111010010",
    "1111001111110110",
    "1111011100010111",
    "1111100111110111",
    "1111110110100010",
    "1111110101001000",
    "1111011100000100",
    "1111000010101011",
    "1110101110110101",
    "1110100101011000",
    "1110101000010011",
    "1110110100101110",
    "1111000100011101",
    "1111010001110000",
    "1111011001000010",
    "1111011011001100",
    "1111011101111011",
    "1111100111111001",
    "1111111100111111",
    "1111100011010101",
    "1110111111001010",
    "1110011110101001",
    "1110001000111110",
    "1110000010000011",
    "1110001000101000",
    "1110010111000011",
    "1110100111010000",
    "1110110100101100",
    "1110111101011100",
    "1111000001110100",
    "1111000010100010",
    "1111000000101100",
    "1110111101001111",
    "1110111000011000",
    "1110110010101011",
    "1110101101010110",
    "1110101001110010",
    "1110101001101011",
    "1110101111011110",
    "1110111101110000",
    "1111010101011111",
    "1111110100110010",
    "1111101000100010",
    "1111000111101101",
    "1110101101100100",
    "1110011101010001",
    "1110010111010000",
    "1110011001001100",
    "1110011111001000",
    "1110100101000000",
    "1110101000001100",
    "1110101000011000",
    "1110100110110100",
    "1110100110000011",
    "1110101010101101",
    "1110111001101011",
    "1111010100101001",
    "1111111001100010",
    "1111011101001100",
    "1110110111000011",
    "1110011010100010",
    "1110001100000010",
    "1110001011110000",
    "1110010101010011",
    "1110100010101110",
    "1110101110101001",
    "1110110110000000",
    "1110111001100010",
    "1110111101000101",
    "1111000101010000",
    "1111010100110100",
    "1111101010100101",
    "1111111110001100",
    "1111101011010001",
    "1111100001001111",
    "1111100001110011",
    "1111101010010000",
    "1111110101010000",
    "1111111101100010",
    "1111111111101001",
    "1111111010011100",
    "1111101110110100",
    "1111011110111101",
    "1111001110000000",
    "1110111110101101",
    "1110110010011111",
    "1110101001110100",
    "1110100100001101",
    "1110100000111110",
    "1110011111101110",
    "1110100000001101",
    "1110100010001101",
    "1110100101100000",
    "1110101001110000",
    "1110101110110110",
    "1110110100101111",
    "1110111100001001",
    "1111000111101111",
    "1111011010110100",
    "1111110110010100",
    "1111100111101111",
    "1111000100100111",
    "1110100110111100",
    "1110010100101001",
    "1110010001000101",
    "1110011011010100",
    "1110101110000010",
    "1111000010100100",
    "1111010010101001",
    "1111011100000010",
    "1111100010111000",
    "1111101101010001",
    "1111111111100101",
    "1111100101010111",
    "1111000101110100",
    "1110101000011011",
    "1110010011101110",
    "1110001100001110",
    "1110010001001111",
    "1110011101101000",
    "1110101011101010",
    "1110111000001001",
    "1111000100000001",
    "1111010010011001",
    "1111100101011000",
    "1111111101000110",
    "1111101000111011",
    "1111010001010010",
    "1110111111111111",
    "1110110110110010",
    "1110110100100111",
    "1110110101111110",
    "1110110111000100",
    "1110110110000001",
    "1110110011111000",
    "1110110100011000",
    "1110111011101010",
    "1111001011110010",
    "1111100011100010",
    "1111111110101100",
    "1111101000011011",
    "1111010110101111",
    "1111001110111011",
    "1111010001001000",
    "1111011011101111",
    "1111101100110101",
    "1111111101001000",
    "1111100100010010",
    "1111001011010001",
    "1110110101011011",
    "1110100101110001",
    "1110011110010001",
    "1110011111100011",
    "1110101000011010",
    "1110110110010110",
    "1111000111011010",
    "1111011010110000",
    "1111110000010001",
    "1111111000011111",
    "1111100001010101",
    "1111001100111000",
    "1110111101110101",
    "1110110110100100",
    "1110110111110001",
    "1111000000001100",
    "1111001101110011",
    "1111011110111101",
    "1111110011001111",
    "1111110101001101",
    "1111011010101000",
    "1110111110010100",
    "1110100011001000",
    "1110001101001100",
    "1110000000011001",
    "1101111110101101",
    "1110000111100010",
    "1110011000001000",
    "1110101100101010",
    "1111000001101001",
    "1111010100111011",
    "1111100110100110",
    "1111111000000010",
    "1111110101100101",
    "1111100010100111",
    "1111010000110011",
    "1111000011000000",
    "1110111011111100",
    "1110111100111000",
    "1111000100110011",
    "1111010000011100",
    "1111011011110101",
    "1111100011010111",
    "1111100100110011",
    "1111011111010111",
    "1111010011110100",
    "1111000100100111",
    "1110110101011000",
    "1110101001110010",
    "1110100100011100",
    "1110100110001001",
    "1110101101101000",
    "1110111000000110",
    "1111000010000000",
    "1111001000011010",
    "1111001010000110",
    "1111001000000001",
    "1111000100101001",
    "1111000011010011",
    "1111001000101100",
    "1111011000110100",
    "1111110100001010",
    "1111101000100001",
    "1111000100000011",
    "1110100110001110",
    "1110010101000000",
    "1110010011001111",
    "1110011111010110",
    "1110110011110011",
    "1111001010010011",
    "1111011101100110",
    "1111101010111001",
    "1111110010010010",
    "1111110101101110",
    "1111111001000110",
    "1111111111001110",
    "1111110001011111",
    "1111011110111010",
    "1111001011010110",
    "1110111100001110",
    "1110110110100111",
    "1110111101110101",
    "1111010010000101",
    "1111110000010101",
    "1111101100101001",
    "1111001011011000",
    "1110110001100010",
    "1110100010100010",
    "1110011110101011",
    "1110100011010101",
    "1110101100011110",
    "1110110101111100",
    "1110111110011110",
    "1111001001011001",
    "1111011011011001",
    "1111110110111100",
    "1111100101010111",
    "1110111111100011",
    "1110011111001010",
    "1110001010101101",
    "1110000110000001",
    "1110001111010111",
    "1110100000100001",
    "1110110010010000",
    "1110111110010111",
    "1111000011101110",
    "1111000111010011",
    "1111001111011110",
    "1111100000100100",
    "1111111010010000",
    "1111101001010100",
    "1111010001111000",
    "1111000101111110",
    "1111001001000100",
    "1111011000111111",
    "1111101111011010",
    "1111111010010110",
    "1111101001001111",
    "1111011110101101",
    "1111011001011110",
    "1111010111101100",
    "1111010111001011",
    "1111010110101100",
    "1111010110111100",
    "1111011001101010",
    "1111100000110001",
    "1111101101110001",
    "1111111111110100",
    "1111101010001010",
    "1111010011101001",
    "1110111110010111",
    "1110101100001100",
    "1110011110111111",
    "1110011000011010",
    "1110011001101000",
    "1110100011010101",
    "1110110101011111",
    "1111001110101101",
    "1111101100010010",
    "1111110101001101",
    "1111011001010101",
    "1111000010100001",
    "1110110010000000",
    "1110100111110010",
    "1110100011000001",
    "1110100010100010",
    "1110100101001000",
    "1110101001110100",
    "1110101111101110",
    "1110110110000001",
    "1110111011100000",
    "1110111110111011",
    "1110111111110000",
    "1110111110010001",
    "1110111011010011",
    "1110110111011011",
    "1110110010111101",
    "1110101110000101",
    "1110101001001011",
    "1110100100101100",
    "1110100001011100",
    "1110100000100111",
    "1110100011101110",
    "1110101100000010",
    "1110111010010001",
    "1111001101101110",
    "1111100100100000",
    "1111111100000001",
    "1111101101110100",
    "1111011010011000",
    "1111001010001011",
    "1110111101011100",
    "1110110100001101",
    "1110101110011100",
    "1110101100011011",
    "1110101110001101",
    "1110110011010010",
    "1110111010010110",
    "1111000001100110",
    "1111000111001101",
    "1111001001110101",
    "1111001001000001",
    "1111000101001000",
    "1110111111010001",
    "1110111000111010",
    "1110110011100010",
    "1110110000000011",
    "1110101110110000",
    "1110110000001111",
    "1110110110001110",
    "1111000010011100",
    "1111010101000101",
    "1111101100000011",
    "1111111100110000",
    "1111101010000111",
    "1111011111100100",
    "1111011110010111",
    "1111100100100010",
    "1111101101100101",
    "1111110100011010",
    "1111110101001110",
    "1111101110111000",
    "1111100010111110",
    "1111010100110111",
    "1111001000010110",
    "1111000000011110",
    "1110111110011110",
    "1111000001110000",
    "1111001000011110",
    "1111010000100001",
    "1111011000001100",
    "1111011110111010",
    "1111100100111001",
    "1111101010111000",
    "1111110010000101",
    "1111111011101010",
    "1111110111100101",
    "1111100111110101",
    "1111010110000110",
    "1111000100010111",
    "1110110100101111",
    "1110101001000110",
    "1110100010001111",
    "1110100000000111",
    "1110100011111110",
    "1110110000011110",
    "1111000110110111",
    "1111100110000000",
    "1111110110010010",
    "1111010100010000",
    "1110111001110100",
    "1110101011010100",
    "1110101010000001",
    "1110110010100001",
    "1110111111010111",
    "1111001011010100",
    "1111010010111110",
    "1111010101101111",
    "1111010101001101",
    "1111010101110001",
    "1111011101011001",
    "1111101111010000",
    "1111110110000111",
    "1111011000010000",
    "1110111110101110",
    "1110101111101011",
    "1110101110000010",
    "1110111000010110",
    "1111001001000100",
    "1111011001101101",
    "1111100101100000",
    "1111101010100011",
    "1111101010000110",
    "1111100110111010",
    "1111100011011100",
    "1111100001001100",
    "1111011111111000",
    "1111011101111010",
    "1111011011010001",
    "1111011010011001",
    "1111011110100011",
    "1111101001110011",
    "1111111011101111",
    "1111101110111110",
    "1111011011010001",
    "1111001101100011",
    "1111000111110100",
    "1111001000011000",
    "1111001011101101",
    "1111001110011111",
    "1111001110101011",
    "1111001100000101",
    "1111001000000110",
    "1111000101010011",
    "1111000111101100",
    "1111010010010000",
    "1111100101010011",
    "1111111110010100",
    "1111100111101011",
    "1111010010010111",
    "1111000110010000",
    "1111000101101001",
    "1111001111111111",
    "1111100010011001",
    "1111111000101100",
    "1111110001101110",
    "1111100000110001",
    "1111010110101010",
    "1111010100001000",
    "1111011000101000",
    "1111100011001101",
    "1111110010101011",
    "1111111010010101",
    "1111100101101010",
    "1111010001100010",
    "1111000000101100",
    "1110110101101111",
    "1110110001111110",
    "1110110101000110",
    "1110111101010001",
    "1111001000000110",
    "1111010011000101",
    "1111011011111101",
    "1111100001010100",
    "1111100010110011",
    "1111100001001000",
    "1111011101101101",
    "1111011001111101",
    "1111010110101100",
    "1111010100010010",
    "1111010010111000",
    "1111010010111011",
    "1111010101011101",
    "1111011011011001",
    "1111100100110110",
    "1111110000111000",
    "1111111101100101",
    "1111110111001000",
    "1111101111000100",
    "1111101011000100",
    "1111101010101011",
    "1111101100010111",
    "1111101110011001",
    "1111101111010111",
    "1111101111000001",
    "1111101110010100",
    "1111101111001111",
    "1111110100000000",
    "1111111110010010",
    "1111110001101010",
    "1111011101100100",
    "1111001000100011",
    "1110110110010101",
    "1110101010010011",
    "1110100110011011",
    "1110101010110101",
    "1110110101110100",
    "1111000100010010",
    "1111010010101111",
    "1111011110100001",
    "1111100110010011",
    "1111101011000110",
    "1111101111110111",
    "1111110111110110",
    "1111111011001000",
    "1111101001110111",
    "1111010111010110",
    "1111000111101000",
    "1110111110011111",
    "1110111110001010",
    "1111000111010000",
    "1111011000111010",
    "1111110001001111",
    "1111110010101001",
    "1111010110000011",
    "1110111100011110",
    "1110101001011101",
    "1110011111100110",
    "1110100000010100",
    "1110101100100000",
    "1111000100100101",
    "1111100111011000",
    "1111101110101001",
    "1111000011101010",
    "1110011110111011",
    "1110000110101111",
    "1101111110100011",
    "1110000110000001",
    "1110011000110100",
    "1110110000100001",
    "1111001000100010",
    "1111100000000010",
    "1111111000010101",
    "1111101101011111",
    "1111010010101100",
    "1110111010110100",
    "1110101010101010",
    "1110100110101101",
    "1110110000100100",
    "1111000101001101",
    "1111011110010100",
    "1111110101000101",
    "1111111011110000",
    "1111110101110101",
    "1111110111100001",
    "1111111101101000",
    "1111111011011111",
    "1111110110101011",
    "1111110101100011",
    "1111111001101100",
    "1111111100000000",
    "1111101100000101",
    "1111011000001011",
    "1111000011001010",
    "1110110000010111",
    "1110100010111110",
    "1110011100111101",
    "1110011101111000",
    "1110100011001010",
    "1110101001011000",
    "1110101101100110",
    "1110101110010111",
    "1110101011111000",
    "1110101001011000",
    "1110101100111010",
    "1110111011100000",
    "1111010110010010",
    "1111111001101100",
    "1111100001100001",
    "1111000011001010",
    "1110110001000101",
    "1110101101011110",
    "1110110101010101",
    "1111000010110110",
    "1111010000100001",
    "1111011010111101",
    "1111100011010000",
    "1111101101100001",
    "1111111100111110",
    "1111101101101111",
    "1111010110010101",
    "1111000011101100",
    "1110111100100000",
    "1111000100111100",
    "1111011100110000",
    "1111111110000010",
    "1111100000000010",
    "1111000101011101",
    "1110110110011101",
    "1110110010101011",
    "1110110111100000",
    "1111000011000011",
    "1111010100010000",
    "1111101010011001",
    "1111111011001101",
    "1111011110110000",
    "1111000011100010",
    "1110101101100001",
    "1110100000011010",
    "1110011101011100",
    "1110100010010000",
    "1110101010110100",
    "1110110011010011",
    "1110111010001011",
    "1111000000100001",
    "1111001000100111",
    "1111010100011100",
    "1111100100110110",
    "1111111000101000",
    "1111110010111111",
    "1111100001010000",
    "1111010101000001",
    "1111001111111101",
    "1111010010101100",
    "1111011101010010",
    "1111101111001100",
    "1111111000111101",
    "1111011101111010",
    "1111000100000000",
    "1110110000011010",
    "1110101000000001",
    "1110101101111111",
    "1111000010001101",
    "1111100000111110",
    "1111111011111111",
    "1111011011110000",
    "1111000011110100",
    "1110110110110111",
    "1110110100100010",
    "1110111010000111",
    "1111000011111100",
    "1111001110100100",
    "1111010111101100",
    "1111011110010110",
    "1111100010101011",
    "1111100101000001",
    "1111100101110110",
    "1111100110000100",
    "1111101000000010",
    "1111101101111110",
    "1111111000101100",
    "1111111001100011",
    "1111101101000111",
    "1111100111100010",
    "1111101101111011",
    "1111111101100111",
    "1111011110010100",
    "1110111011100011",
    "1110011101111111",
    "1110001100100011",
    "1110001010000111",
    "1110010101001000",
    "1110101000101100",
    "1111000000001101",
    "1111011010110101",
    "1111111001111010",
    "1111100001111001",
    "1110111010001001",
    "1110010011100111",
    "1101110100110111",
    "1101100100001010",
    "1101100100111100",
    "1101110101001000",
    "1110001110000101",
    "1110101000010011",
    "1110111101100100",
    "1111001011000111",
    "1111010001100111",
    "1111010101010011",
    "1111011100101000",
    "1111101100010110",
    "1111111011001111",
    "1111011101111101",
    "1111000001111001",
    "1110101100111000",
    "1110100010010100",
    "1110100010011001",
    "1110101001110101",
    "1110110100010111",
    "1110111110010111",
    "1111000101100101",
    "1111001001011110",
    "1111001010100101",
    "1111001010111000",
    "1111001110011001",
    "1111011000110111",
    "1111101011101000",
    "1111111010101101",
    "1111011110011001",
    "1111000100100101",
    "1110110001110001",
    "1110101000010001",
    "1110100111001110",
    "1110101011100001",
    "1110110001111101",
    "1110111000001110",
    "1110111101110000",
    "1111000011011111",
    "1111001010011011",
    "1111010010010000",
    "1111011000110100",
    "1111011010010011",
    "1111010011100010",
    "1111000100010011",
    "1110101111100011",
    "1110011010010110",
    "1110001010010011",
    "1110000010111110",
    "1110000100111001",
    "1110001110000000",
    "1110011010111111",
    "1110101000110101",
    "1110110101011011",
    "1111000001000000",
    "1111001111101011",
    "1111100110000100",
    "1111111010001001",
    "1111010011011100",
    "1110101100100000",
    "1110001101010111",
    "1101111100011011",
    "1101111100101011",
    "1110001011011011",
    "1110100001011111",
    "1110110111011111",
    "1111001000010011",
    "1111010100011100",
    "1111100001000111",
    "1111110011010101",
    "1111110010101101",
    "1111010011110100",
    "1110110111110010",
    "1110100111110010",
    "1110101011000111",
    "1111000011111100",
    "1111101100111110",
    "1111100100000101",
    "1110111010010001",
    "1110011101100100",
    "1110010000010101",
    "1110010000011001",
    "1110011001101000",
    "1110101000101000",
    "1110111011101111",
    "1111010010001000",
    "1111101010101110",
    "1111111100101001",
    "1111100111000110",
    "1111011000010000",
    "1111010010111011",
    "1111010110110110",
    "1111100000110000",
    "1111101100100111",
    "1111110111001010",
    "1111111111011101",
    "1111111000010011",
    "1111101100101100",
    "1111011011000100",
    "1111000011111100",
    "1110101011110111",
    "1110011001100111",
    "1110010011101010",
    "1110011110001100",
    "1110111001010000",
    "1111100000101100",
    "1111110001111000",
    "1111000101100100",
    "1110100000001010",
    "1110000101010011",
    "1101110110100010",
    "1101110011011010",
    "1101111001110111",
    "1110000111010001",
    "1110011000011110",
    "1110101010010110",
    "1110111010101010",
    "1111001000010001",
    "1111010101001001",
    "1111100101111110",
    "1111111110011100",
    "1111100000110101",
    "1110111011100000",
    "1110011000101111",
    "1101111111110110",
    "1101110101111011",
    "1101111011101000",
    "1110001011110000",
    "1110011110100110",
    "1110101101010111",
    "1110110101001011",
    "1110111001100101",
    "1111000000110011",
    "1111001111010100",
    "1111100110000001",
    "1111111111101000",
    "1111101010000000",
    "1111100001001101",
    "1111101010101000",
    "1111111010101000",
    "1111010110001001",
    "1110110010001101",
    "1110011000011011",
    "1110001110011011",
    "1110010101011111",
    "1110101011110111",
    "1111001101000111",
    "1111110011001111",
    "1111100111010100",
    "1111000110110110",
    "1110101110010001",
    "1110011110111010",
    "1110011000111001",
    "1110011011010001",
    "1110100100000110",
    "1110110000100001",
    "1110111101011110",
    "1111001000011101",
    "1111010000011001",
    "1111010101011011",
    "1111011000101010",
    "1111011100100000",
    "1111100100001000",
    "1111110010001111",
    "1111110111111111",
    "1111011100001001",
    "1110111101110011",
    "1110100001101110",
    "1110001100011110",
    "1110000000110101",
    "1101111110110101",
    "1110000100001010",
    "1110001101000010",
    "1110010101111100",
    "1110011100111000",
    "1110100001001100",
    "1110100011010000",
    "1110100100001000",
    "1110100101100100",
    "1110101010000010",
    "1110110011111011",
    "1111000100011100",
    "1111011011000110",
    "1111110101100110",
    "1111101111011010",
    "1111010111101111",
    "1111000110110001",
    "1110111110010010",
    "1110111110001010",
    "1111000101000101",
    "1111010001100110",
    "1111100010101011",
    "1111110111000110",
    "1111110011001100",
    "1111011111101001",
    "1111010010000110",
    "1111001110000101",
    "1111010101110001",
    "1111101000110011",
    "1111111100000011",
    "1111011110001010",
    "1111000011010111",
    "1110110000011110",
    "1110101000110010",
    "1110101110010010",
    "1111000000111101",
    "1111011110010001",
    "1111111110010010",
    "1111011010110000",
    "1110111100111100",
    "1110101001010001",
    "1110100001110001",
    "1110100101001001",
    "1110101111101000",
    "1110111100001001",
    "1111000111011101",
    "1111010010001101",
    "1111011111010111",
    "1111110001101000",
    "1111110110011000",
    "1111011011000111",
    "1111000000111101",
    "1110101100100110",
    "1110100001010000",
    "1110011110110101",
    "1110100010010101",
    "1110101000110010",
    "1110110001011111",
    "1110111110110101",
    "1111010100010010",
    "1111110010111111",
    "1111100111011110",
    "1111000000111101",
    "1110100001001101",
    "1110001111010110",
    "1110001111000000",
    "1110011111010100",
    "1110111011001010",
    "1111011011011001",
    "1111111001011110",
    "1111101110110001",
    "1111011111001100",
    "1111010111111111",
    "1111011000100011",
    "1111011111111111",
    "1111101100111101",
    "1111111101110000",
    "1111101111100011",
    "1111011101001111",
    "1111001101001100",
    "1111000000111001",
    "1110111000111111",
    "1110110101001001",
    "1110110100110110",
    "1110110111101010",
    "1110111101011011",
    "1111000101100101",
    "1111001111001111",
    "1111011001001110",
    "1111100010011101",
    "1111101010010001",
    "1111110000000011",
    "1111110100010000",
    "1111111010101110",
    "1111110111100010",
    "1111100000100110",
    "1111000010100111",
    "1110100100010000",
    "1110001101110101",
    "1110000101101010",
    "1110001110101110",
    "1110100110000100",
    "1111000011100100",
    "1111011110010100",
    "1111101111011011",
    "1111110110001010",
    "1111111000011011",
    "1111111101000000",
    "1111110111110010",
    "1111100101101111",
    "1111010001101110",
    "1111000010001000",
    "1110111100001110",
    "1111000010001101",
    "1111010000101011",
    "1111100000111011",
    "1111101101001010",
    "1111110010100010",
    "1111110010010111",
    "1111110000000101",
    "1111101110011010",
    "1111110000001001",
    "1111111000100111",
    "1111110110001111",
    "1111011100110111",
    "1110111110000111",
    "1110011111011010",
    "1110000110010011",
    "1101110111011000",
    "1101110101100010",
    "1110000000000111",
    "1110010010101011",
    "1110100111001011",
    "1110110111110111",
    "1111000001100100",
    "1111000100010101",
    "1111000010010101",
    "1111000001000011",
    "1111000111000001",
    "1111010111010110",
    "1111110001000000",
    "1111110001001000",
    "1111010110001001",
    "1111000011100010",
    "1110111100000100",
    "1110111111000100",
    "1111001000101010",
    "1111010100010101",
    "1111011110011110",
    "1111100101100111",
    "1111101011011100",
    "1111110010100101",
    "1111111100100100",
    "1111110110111110",
    "1111101010100010",
    "1111100000110011",
    "1111011011000110",
    "1111011000111010",
    "1111010111101100",
    "1111010011101001",
    "1111001001100011",
    "1110111000110101",
    "1110100100000110",
    "1110001111111011",
    "1110000000100001",
    "1101111000101000",
    "1101111001000110",
    "1110000001000010",
    "1110001111110110",
    "1110100110001011",
    "1111000011111011",
    "1111100111011101",
    "1111110010100110",
    "1111001111110110",
    "1110110101111011",
    "1110101001001011",
    "1110101010100011",
    "1110110110111001",
    "1111001001111101",
    "1111100000011111",
    "1111111000000000",
    "1111110000111000",
    "1111011011111111",
    "1111001011011110",
    "1111000001001101",
    "1110111111000010",
    "1111000101110110",
    "1111010100001011",
    "1111100111000011",
    "1111111010011011",
    "1111110101010000",
    "1111101010001111",
    "1111100100111011",
    "1111100100010101",
    "1111100110101011",
    "1111101010101111",
    "1111110000010000",
    "1111110111011111",
    "1111111111010110",
    "1111110100111010",
    "1111101010101100",
    "1111100010011100",
    "1111011101010100",
    "1111011011100011",
    "1111011100110011",
    "1111100000100100",
    "1111100110011010",
    "1111101101110011",
    "1111110110100000",
    "1111111111110110",
    "1111110110001011",
    "1111101101101111",
    "1111101000000000",
    "1111100101110111",
    "1111100110111001",
    "1111101000110000",
    "1111101000000001",
    "1111100001100001",
    "1111010011110110",
    "1111000000001101",
    "1110101010100000",
    "1110010111111010",
    "1110001100110010",
    "1110001011001110",
    "1110010010100100",
    "1110100000101001",
    "1110110100111100",
    "1111010000001010",
    "1111110010000010",
    "1111100111010100",
    "1111000000100011",
    "1110011111100001",
    "1110001001001011",
    "1110000000101100",
    "1110000101001011",
    "1110010001100010",
    "1110011111111101",
    "1110101011100011",
    "1110110010001011",
    "1110110100110100",
    "1110110101100000",
    "1110110110010010",
    "1110111000100111",
    "1110111100010100",
    "1111000001110011",
    "1111001011011110",
    "1111011011101111",
    "1111110011101100",
    "1111101101110100",
    "1111001101000101",
    "1110110000000010",
    "1110011100101010",
    "1110010110011101",
    "1110011100001001",
    "1110101000111010",
    "1110110111001110",
    "1111000010011001",
    "1111001000010000",
    "1111001000111111",
    "1111000110001110",
    "1111000010010101",
    "1110111111001100",
    "1110111101000111",
    "1110111011110101",
    "1110111010110111",
    "1110111001111101",
    "1110111001101101",
    "1110111010111010",
    "1110111101111000",
    "1111000001111110",
    "1111000101110010",
    "1111001000000100",
    "1111001000110111",
    "1111001001110000",
    "1111001101110000",
    "1111010111110010",
    "1111101001000101",
    "1111111111100110",
    "1111100101101010",
    "1111001101010010",
    "1110111010000111",
    "1110101110001100",
    "1110101001110000",
    "1110101011101010",
    "1110110001110000",
    "1110111010000111",
    "1111000011011101",
    "1111001101001001",
    "1111011000001100",
    "1111100110111011",
    "1111111010100011",
    "1111101101110110",
    "1111010101101010",
    "1111000001100110",
    "1110110101100111",
    "1110110100001101",
    "1110111101011100",
    "1111001110110001",
    "1111100100011101",
    "1111111010111010",
    "1111110000110000",
    "1111100000011100",
    "1111010101010101",
    "1111010000001010",
    "1111010000101110",
    "1111010110100000",
    "1111100000110011",
    "1111101110010110",
    "1111111101100110",
    "1111110011010001",
    "1111100110011011",
    "1111011101111011",
    "1111011011101000",
    "1111100000100100",
    "1111101100101001",
    "1111111110010111",
    "1111101100110110",
    "1111011000011110",
    "1111000111101000",
    "1110111100010100",
    "1110110110111011",
    "1110110110000001",
    "1110110111100000",
    "1110111001101010",
    "1110111011100000",
    "1110111101000100",
    "1110111110101101",
    "1111000000110000",
    "1111000011010111",
    "1111000110001101",
    "1111001001001011",
    "1111001110001111",
    "1111011000110000",
    "1111101010101101",
    "1111111100010111",
    "1111100000010111",
    "1111000111010011",
    "1110110111001000",
    "1110110100000011",
    "1110111110010100",
    "1111010001001000",
    "1111100101101100",
    "1111110101010111",
    "1111111100111011",
    "1111111111011100",
    "1111111101011000",
    "1111110100111110",
    "1111100101100010",
    "1111010001111110",
    "1110111111110110",
    "1110110100110001",
    "1110110110001011",
    "1111000111000100",
    "1111100101100101",
    "1111110011011001",
    "1111001010111101",
    "1110101000000011",
    "1110001111011010",
    "1110000100010000",
    "1110000110101100",
    "1110010010110011",
    "1110100101100010",
    "1110111110001001",
    "1111011100000001",
    "1111111110100000",
    "1111011101001111",
    "1110111100110000",
    "1110100100110001",
    "1110011000111100",
    "1110011010100011",
    "1110100110101101",
    "1110111000011011",
    "1111001010101011",
    "1111011001000010",
    "1111100010010010",
    "1111101000100110",
    "1111101111111110",
    "1111111100000110",
    "1111110010101001",
    "1111011111111011",
    "1111010000101110",
    "1111001001100011",
    "1111001100101101",
    "1111011000101000",
    "1111101001000100",
    "1111111001100001",
    "1111111000110000",
    "1111101110000100",
    "1111100101001110",
    "1111011101010010",
    "1111010101100111",
    "1111001110010110",
    "1111001000101000",
    "1111000101111110",
    "1111000111100111",
    "1111001110000000",
    "1111011001011101",
    "1111101011000000",
    "1111111100101001",
    "1111011110100100",
    "1110111101110101",
    "1110011111011111",
    "1110001001000100",
    "1101111110100110",
    "1110000001001100",
    "1110001101110101",
    "1110011110111111",
    "1110101111001100",
    "1110111010110100",
    "1111000001000000",
    "1111000010111101",
    "1111000010101001",
    "1111000010000010",
    "1111000010011100",
    "1111000100101110",
    "1111001001011011",
    "1111010000010101",
    "1111011000000110",
    "1111011110010100",
    "1111100000010010",
    "1111011011101101",
    "1111001111100100",
    "1110111101011001",
    "1110101001100111",
    "1110011001111100",
    "1110010011010000",
    "1110010111011111",
    "1110100101001110",
    "1110111010000110",
    "1111010100010101",
    "1111110010001111",
    "1111101110001111",
    "1111010000000000",
    "1110110110101100",
    "1110100101100101",
    "1110011110110000",
    "1110100010001011",
    "1110101100100110",
    "1110111001001011",
    "1111000011011100",
    "1111001000110111",
    "1111001011001111",
    "1111001111111010",
    "1111011011101011",
    "1111110000101001",
    "1111110011010100",
    "1111010110100101",
    "1110111111111101",
    "1110110100110111",
    "1110110111010101",
    "1111000100011101",
    "1111010111000001",
    "1111101010001010",
    "1111111011001110",
    "1111110101111111",
    "1111101000111010",
    "1111011101001111",
    "1111010010110011",
    "1111001010010001",
    "1111000101011111",
    "1111000110001101",
    "1111001101110011",
    "1111011100110101",
    "1111110010010010",
    "1111110100000010",
    "1111011001000111",
    "1110111111111111",
    "1110101011011001",
    "1110011101101000",
    "1110011000001100",
    "1110011010111111",
    "1110100100011000",
    "1110110001101100",
    "1111000000000010",
    "1111001110010110",
    "1111011110001101",
    "1111110001110100",
    "1111110101011000",
    "1111011000010110",
    "1110111010100000",
    "1110100000110001",
    "1110010000000011",
    "1110001011000111",
    "1110010001100100",
    "1110100010100100",
    "1110111101101000",
    "1111100000111001",
    "1111110110111011",
    "1111001110110011",
    "1110101100101110",
    "1110010101110100",
    "1110001101100110",
    "1110010100110110",
    "1110100111101000",
    "1111000001001101",
    "1111011111101000",
    "1111111101111110",
    "1111011000011101",
    "1110110001111110",
    "1110001111000111",
    "1101110100100010",
    "1101100110011000",
    "1101100111000011",
    "1101110100000101",
    "1110000111110010",
    "1110011110010110",
    "1110110110110100",
    "1111010010011100",
    "1111110010110011",
    "1111101001000101",
    "1111000101010000",
    "1110100111010101",
    "1110010101110110",
    "1110010100001011",
    "1110100000010010",
    "1110110100011111",
    "1111001001101111",
    "1111011010010011",
    "1111100101001000",
    "1111101101000011",
    "1111110110011101",
    "1111111011000011",
    "1111100111110011",
    "1111010011011111",
    "1111000010110110",
    "1110111001110010",
    "1110111001110000",
    "1111000000110001",
    "1111001010111000",
    "1111010100100101",
    "1111011101011110",
    "1111101000010000",
    "1111110111111100",
    "1111110010100100",
    "1111011001011101",
    "1111000001010101",
    "1110101111110110",
    "1110101001000100",
    "1110101101111011",
    "1110111011100110",
    "1111001100111000",
    "1111011100101101",
    "1111101000001001",
    "1111101110110110",
    "1111110010000011",
    "1111110011101000",
    "1111110101011011",
    "1111111000101111",
    "1111111110001011",
    "1111111010100001",
    "1111110010101001",
    "1111101100010111",
    "1111101010011010",
    "1111101110111111",
    "1111111011010101",
    "1111110001000110",
    "1111011001100010",
    "1111000010110110",
    "1110110010001000",
    "1110101010101010",
    "1110101101000100",
    "1110110111100011",
    "1111000110101000",
    "1111010110010011",
    "1111100011010111",
    "1111101101011011",
    "1111110111110001",
    "1111111001000101",
    "1111100010110100",
    "1111000110110001",
    "1110101001110101",
    "1110010010100010",
    "1110000110111111",
    "1110001011001110",
    "1110011110101001",
    "1110111011111010",
    "1111011011011011",
    "1111110101110111",
    "1111111001010101",
    "1111110011100011",
    "1111110111110011",
    "1111111100011110",
    "1111101100110001",
    "1111011011111000",
    "1111001011110010",
    "1110111101100011",
    "1110110001111000",
    "1110101001110100",
    "1110100110011011",
    "1110101000100111",
    "1110110000010101",
    "1110111100111100",
    "1111001101011110",
    "1111100000111011",
    "1111110101111010",
    "1111110101000001",
    "1111100001010000",
    "1111001111101001",
    "1111000000101100",
    "1110110100111011",
    "1110101101000111",
    "1110101010001110",
    "1110101101101000",
    "1110111000110010",
    "1111001100001110",
    "1111100110111000",
    "1111111001111101",
    "1111011010001001",
    "1110111101001111",
    "1110100110000000",
    "1110010110000000",
    "1110001101100100",
    "1110001011111111",
    "1110001111111101",
    "1110010111110101",
    "1110100001111110",
    "1110101100101101",
    "1110110110001101",
    "1110111110000000",
    "1111000110101010",
    "1111010011101110",
    "1111100110111000",
    "1111111110111101",
    "1111101000101001",
    "1111010101110111",
    "1111001110101110",
    "1111011001010000",
    "1111110111000101",
    "1111011100010100",
    "1110101001111101",
    "1101111100111101",
    "1101011110011110",
    "1101010010110110",
    "1101011010001001",
    "1101101111010010",
    "1110001010001100",
    "1110100011111100",
    "1110111000010011",
    "1111000110000011",
    "1111010000011111",
    "1111011101101000",
    "1111110010010110",
    "1111110000000101",
    "1111001101010001",
    "1110101100010111",
    "1110010101000110",
    "1110001101100011",
    "1110010111100011",
    "1110101110011110",
    "1111001010001011",
    "1111100010111011",
    "1111110011100011",
    "1111111010110110",
    "1111111010011111",
    "1111110101010000",
    "1111101110101100",
    "1111101001000001",
    "1111100100010010",
    "1111011111100011",
    "1111011010100110",
    "1111011000010000",
    "1111011100101011",
    "1111101010001100",
    "1111111111101101",
    "1111100111101011",
    "1111010010110011",
    "1111000111001101",
    "1111000111011011",
    "1111010001011110",
    "1111011111101011",
    "1111101100010100",
    "1111110100010001",
    "1111111000111011",
    "1111111110110101",
    "1111110110000000",
    "1111100100010101",
    "1111001110001101",
    "1110111000101000",
    "1110101000111111",
    "1110100011001111",
    "1110101000101100",
    "1110110111010110",
    "1111001011100011",
    "1111100001110011",
    "1111111000000101",
    "1111110010110101",
    "1111100000111001",
    "1111010100010000",
    "1111001101111011",
    "1111001101001111",
    "1111010000000111",
    "1111010011100110",
    "1111010101001001",
    "1111010011101110",
    "1111001111110110",
    "1111001011011101",
    "1111001001000111",
    "1111001010111010",
    "1111010001000111",
    "1111011010000001",
    "1111100010101111",
    "1111101000111100",
    "1111101011110110",
    "1111101100101010",
    "1111101110001001",
    "1111110011001001",
    "1111111101011110",
    "1111110010110010",
    "1111011111110000",
    "1111001100101010",
    "1110111100011110",
    "1110110001000010",
    "1110101010010011",
    "1110100110111001",
    "1110100100111011",
    "1110100010100010",
    "1110011110111101",
    "1110011010011101",
    "1110010110011000",
    "1110010100000000",
    "1110010101000000",
    "1110011011101111",
    "1110101010001100",
    "1111000000111001",
    "1111011101111010",
    "1111111101000101",
    "1111100110011101",
    "1111010001010101",
    "1111000110010011",
    "1111000101000000",
    "1111001010101011",
    "1111010011011100",
    "1111011011101011",
    "1111100001001101",
    "1111100011000001",
    "1111100001011110",
    "1111011101101000",
    "1111011000101010",
    "1111010011011100",
    "1111001110110001",
    "1111001011001111",
    "1111001001100010",
    "1111001010110000",
    "1111010000010001",
    "1111011010011101",
    "1111101000011100",
    "1111111000010010",
    "1111110111110001",
    "1111101000100001",
    "1111011001100101",
    "1111001001100011",
    "1110110110110001",
    "1110100000110001",
    "1110001001001001",
    "1101110011000110",
    "1101100010101111",
    "1101011011000100",
    "1101011101001100",
    "1101100111111111",
    "1101111000100101",
    "1110001011001100",
    "1110011100111000",
    "1110101011111101",
    "1110110111111111",
    "1111000011000000",
    "1111010001000111",
    "1111100101010011",
    "1111111111110000",
    "1111100010101011",
    "1111000111101111",
    "1110110101000000",
    "1110101110100001",
    "1110110101010000",
    "1111000101010000",
    "1111011000000100",
    "1111100111101101",
    "1111101111110111",
    "1111101111101110",
    "1111101000111100",
    "1111011110011100",
    "1111010100000001",
    "1111001100101110",
    "1111001011100000",
    "1111010011111110",
    "1111100111110100",
    "1111111010100010",
    "1111010111100111",
    "1110110110010110",
    "1110011101100100",
    "1110010010001000",
    "1110010101000001",
    "1110100001111110",
    "1110110010000101",
    "1111000000110001",
    "1111001110001101",
    "1111011101101011",
    "1111110010001111",
    "1111110100000011",
    "1111011000011110",
    "1111000000011001",
    "1110110001100001",
    "1110101111010001",
    "1110111001110100",
    "1111001111010110",
    "1111101100000110",
    "1111110100100011",
    "1111010110101100",
    "1110111101100110",
    "1110101011111101",
    "1110100011001000",
    "1110100011001010",
    "1110101010000001",
    "1110110100000110",
    "1110111101110011",
    "1111000100101001",
    "1111001001101010",
    "1111010000100100",
    "1111011100111100",
    "1111110000110101",
    "1111110101001010",
    "1111011010001110",
    "1111000100111011",
    "1110111011100011",
    "1111000010000011",
    "1111011000100000",
    "1111111011011110",
    "1111011011001001",
    "1110110010110011",
    "1110010010000010",
    "1101111101101101",
    "1101111000001011",
    "1110000001001101",
    "1110010111010000",
    "1110110111111111",
    "1111100000000111",
    "1111110100100000",
    "1111001010101101",
    "1110100111100111",
    "1110001111101001",
    "1110000101011111",
    "1110001001100000",
    "1110011001111010",
    "1110110011000011",
    "1111010000011111",
    "1111101101110101",
    "1111111000100010",
    "1111100101001001",
    "1111011000111111",
    "1111010011011010",
    "1111010010101110",
    "1111010101011000",
    "1111011010011011",
    "1111100001100001",
    "1111101010010110",
    "1111110100011101",
    "1111111111010000",
    "1111110101111000",
    "1111101011110101",
    "1111100011100111",
    "1111011110110011",
    "1111011111001100",
    "1111100110000110",
    "1111110011110011",
    "1111111000100110",
    "1111100001001111",
    "1111001000111010",
    "1110110011001000",
    "1110100011010101",
    "1110011100000111",
    "1110011110011001",
    "1110101001010110",
    "1110111011000001",
    "1111010000110011",
    "1111101000001100",
    "1111111111000000",
    "1111101100011001",
    "1111011001011101",
    "1111000101101010",
    "1110101111001101",
    "1110010110010011",
    "1101111110000101",
    "1101101011101000",
    "1101100011101111",
    "1101101001010101",
    "1101111011100110",
    "1110010101011010",
    "1110101111110001",
    "1111000100011010",
    "1111010001001100",
    "1111011010010100",
    "1111100101111011",
    "1111111000010000",
    "1111101110000100",
    "1111010001110000",
    "1110111001110101",
    "1110101100111111",
    "1110101111001100",
    "1110111111110101",
    "1111011011110000",
    "1111111110110011",
    "1111011011110101",
    "1110111000001011",
    "1110011010000100",
    "1110000101100100",
    "1101111101000100",
    "1110000000101110",
    "1110001101101101",
    "1110011110011111",
    "1110101101010111",
    "1110110110000100",
    "1110110110111111",
    "1110110001010010",
    "1110100111111111",
    "1110011111010001",
    "1110011010100011",
    "1110011011110010",
    "1110100100011000",
    "1110110101000000",
    "1111001100100000",
    "1111101000010011",
    "1111111011001010",
    "1111100010000000",
    "1111001111111011",
    "1111000111001001",
    "1111000111001101",
    "1111001101001010",
    "1111010110000011",
    "1111100001000010",
    "1111101111000011",
    "1111111110111111",
    "1111101010000100",
    "1111010101100101",
    "1111000110100000",
    "1111000001111001",
    "1111001011010011",
    "1111100010001011",
    "1111111101110101",
    "1111011011011110",
    "1110111101110011",
    "1110101001111111",
    "1110100001111011",
    "1110100100110100",
    "1110101111101100",
    "1110111111101000",
    "1111010011100001",
    "1111101011010110",
    "1111111000110110",
    "1111011001111111",
    "1110111010011011",
    "1110011101010111",
    "1110000110001011",
    "1101110111001011",
    "1101110000110001",
    "1101110001111001",
    "1101111001000010",
    "1110000101010010",
    "1110011000000110",
    "1110110100000001",
    "1111011001101011",
    "1111111001011100",
    "1111001011010100",
    "1110100011101001",
    "1110001000110100",
    "1101111110010110",
    "1110000100010011",
    "1110010111111111",
    "1110110101011101",
    "1111011000001100",
    "1111111011111110",
    "1111100010111110",
    "1111001000101111",
    "1110111000110010",
    "1110110100111011",
    "1110111110001010",
    "1111010100001000",
    "1111110100001010",
    "1111100110010101",
    "1111000001011001",
    "1110100011001000",
    "1110010000001000",
    "1110001010000111",
    "1110001111011111",
    "1110011100001100",
    "1110101011011110",
    "1110111001111100",
    "1111000111100010",
    "1111010111011010",
    "1111101100110001",
    "1111110110111111",
    "1111010101010000",
    "1110110010011101",
    "1110010100101110",
    "1110000001100100",
    "1101111011111010",
    "1110000010100110",
    "1110010001100100",
    "1110100100010111",
    "1110110111011011",
    "1111001001010110",
    "1111011001101111",
    "1111101000111010",
    "1111111001010000",
    "1111110010011110",
    "1111011001101011",
    "1110111110001001",
    "1110100100010010",
    "1110010001111000",
    "1110001011101000",
    "1110010011101010",
    "1110101000000011",
    "1111000010111110",
    "1111011101010111",
    "1111110000110100",
    "1111111001011111",
    "1111110111001011",
    "1111101100010001",
    "1111011101000100",
    "1111001110010111",
    "1111000011011101",
    "1110111101010001",
    "1110111011000001",
    "1110111010110010",
    "1110111010111000",
    "1110111010101000",
    "1110111010001100",
    "1110111010000010",
    "1110111010101101",
    "1110111100101010",
    "1111000000000010",
    "1111000110011111",
    "1111010011001011",
    "1111101000011101",
    "1111111001110101",
    "1111010111010001",
    "1110110101111011",
    "1110011100000010",
    "1110001110101001",
    "1110001111110000",
    "1110011100001100",
    "1110101101111010",
    "1110111111000010",
    "1111001101101110",
    "1111011100111010",
    "1111110000010101",
    "1111110110010101",
    "1111011000100101",
    "1110111011011001",
    "1110100101000110",
    "1110011010101111",
    "1110011101101101",
    "1110101010100010",
    "1110111011001100",
    "1111001001111001",
    "1111010011000000",
    "1111010110011101",
    "1111010110010011",
    "1111010110011101",
    "1111011100011001",
    "1111101011111100",
    "1111111010011011",
    "1111011001100111",
    "1110110111001000",
    "1110011001010110",
    "1110000101101111",
    "1101111111010010",
    "1110000101100100",
    "1110010101010101",
    "1110101001110100",
    "1110111101101110",
    "1111001101000100",
    "1111010101110110",
    "1111010111111111",
    "1111010101001101",
    "1111001111101110",
    "1111001001010011",
    "1111000010101110",
    "1110111011110010",
    "1110110011101111",
    "1110101010011001",
    "1110100000100100",
    "1110010111111010",
    "1110010010011100",
    "1110010001110011",
    "1110010110101100",
    "1110100000111001",
    "1110110000111000",
    "1111000111010101",
    "1111100011111011",
    "1111111011000100",
    "1111011000111110",
    "1110111001111001",
    "1110100010010010",
    "1110010101111100",
    "1110010101110100",
    "1110011111011110",
    "1110101110101110",
    "1110111111011010",
    "1111001110011100",
    "1111011010111100",
    "1111100111000111",
    "1111110111000111",
    "1111110010001111",
    "1111010101110111",
    "1110111000001110",
    "1110011111100011",
    "1110010001100110",
    "1110010010000110",
    "1110100001001000",
    "1110111011001001",
    "1111011011010100",
    "1111111100100000",
    "1111100101110111",
    "1111001111000100",
    "1111000001001100",
    "1110111101001010",
    "1111000010000011",
    "1111001101111010",
    "1111011110000100",
    "1111101111100101",
    "1111111111101011",
    "1111110001010011",
    "1111100110001011",
    "1111011110011111",
    "1111011001110010",
    "1111010111001011",
    "1111010110001000",
    "1111010110110100",
    "1111011001100000",
    "1111011101110011",
    "1111100010111000",
    "1111100111100001",
    "1111101011001001",
    "1111101110000010",
    "1111110001000000",
    "1111110100110011",
    "1111111001101100",
    "1111111111000011",
    "1111111100101101",
    "1111111011011010",
    "1111111110001000",
    "1111111011001001",
    "1111110001100110",
    "1111100111001011",
    "1111011110101011",
    "1111011010111010",
    "1111011101100110",
    "1111100110100001",
    "1111110011111111",
    "1111111100010001",
    "1111101100000001",
    "1111011011110111",
    "1111001011011011",
    "1110111001110000",
    "1110100110100000",
    "1110010010111101",
    "1110000001101110",
    "1101110110000001",
    "1101110010010000",
    "1101110110101000",
    "1110000001000000",
    "1110001101101001",
    "1110011000100010",
    "1110011111000111",
    "1110100000111001",
    "1110011111011001",
    "1110011111001101",
    "1110100110110100",
    "1110111010000100",
    "1111011000100111",
    "1111111101010100",
    "1111011111100110",
    "1111000101010000",
    "1110111000100010",
    "1110111010000111",
    "1111000101110010",
    "1111010101100010",
    "1111100100010111",
    "1111110000100001",
    "1111111100000011",
    "1111110110101010",
    "1111100111011001",
    "1111010111111001",
    "1111001011101111",
    "1111000110010011",
    "1111001000100010",
    "1111010000011010",
    "1111011001011000",
    "1111011110010111",
    "1111011100110000",
    "1111010101011011",
    "1111001100011001",
    "1111000110011111",
    "1111000110110111",
    "1111001110100100",
    "1111011100101010",
    "1111101110100111",
    "1111111110110111",
    "1111101111001001",
    "1111100100110111",
    "1111100001010101",
    "1111100101000101",
    "1111110001010000",
    "1111111001010010",
    "1111011100000001",
    "1110111010111100",
    "1110011011110111",
    "1110000100100111",
    "1101111001100011",
    "1101111100100110",
    "1110001011110011",
    "1110100001110110",
    "1110111000100101",
    "1111001010111000",
    "1111010110000100",
    "1111011001111100",
    "1111010111100000",
    "1111010000110000",
    "1111001000111001",
    "1111000011111011",
    "1111000101001101",
    "1111001110000101",
    "1111011101000111",
    "1111101110100001",
    "1111111101110000",
    "1111111001100000",
    "1111111010001000",
    "1111111100001100",
    "1111101101001100",
    "1111011110001001",
    "1111010011110001",
    "1111010000100100",
    "1111010100111001",
    "1111011111100100",
    "1111101110100111",
    "1111111111101101",
    "1111101111000001",
    "1111011111001000",
    "1111010001110001",
    "1111001000000100",
    "1111000011001111",
    "1111000100001110",
    "1111001011000111",
    "1111010110100111",
    "1111100100100101",
    "1111110010001100",
    "1111111100010111",
    "1111111111100100",
    "1111111100110011",
    "1111110010000101",
    "1111100010101011",
    "1111010010011100",
    "1111000101101110",
    "1111000000010100",
    "1111000100110001",
    "1111010011011000",
    "1111101001111000",
    "1111111011111100",
    "1111100010110110",
    "1111001110110000",
    "1111000001110100",
    "1110111100010001",
    "1110111100110011",
    "1111000000111101",
    "1111000110000011",
    "1111001001111111",
    "1111001011101000",
    "1111001010110010",
    "1111000111110111",
    "1111000011101100",
    "1110111111010110",
    "1110111011111101",
    "1110111010101111",
    "1110111100100101",
    "1111000010010010",
    "1111001100101110",
    "1111011100011001",
    "1111110001000100",
    "1111110110110001",
    "1111011101111101",
    "1111000111001001",
    "1110110100010111",
    "1110100110110100",
    "1110011110111111",
    "1110011100011001",
    "1110011101101101",
    "1110100000111000",
    "1110100100001000",
    "1110100110000001",
    "1110100101110111",
    "1110100110001011",
    "1110101011101111",
    "1110111010000001",
    "1111010001101011",
    "1111101111010011",
    "1111110011011010",
    "1111011100111000",
    "1111010010010100",
    "1111010100111110",
    "1111100001110011",
    "1111110110000001",
    "1111101111110100",
    "1111010001011001",
    "1110110000010001",
    "1110010000000010",
    "1101110101111001",
    "1101100110010011",
    "1101100101100111",
    "1101110110011011",
    "1110010111010110",
    "1111000011101110",
    "1111110100000011",
    "1111100000001010",
    "1110111111011001",
    "1110101101001010",
    "1110101001011110",
    "1110110001000111",
    "1110111111011010",
    "1111001111111111",
    "1111011111000111",
    "1111101011000010",
    "1111110011101101",
    "1111111001100101",
    "1111111101101011",
    "1111111110110001",
    "1111111010111111",
    "1111110110110100",
    "1111110001101010",
    "1111101000111000",
    "1111011001100000",
    "1111000010100100",
    "1110100110011011",
    "1110001010111100",
    "1101110111010001",
    "1101110000110101",
    "1101111001010000",
    "1110001101000111",
    "1110100101011011",
    "1110111010101101",
    "1111000111001001",
    "1111001010010001",
    "1111001001001001",
    "1111001001110111",
    "1111010001000011",
    "1111011111111011",
    "1111110011010100",
    "1111111001110001",
    "1111101100010111",
    "1111100111001011",
    "1111101000011010",
    "1111101011101111",
    "1111101101001010",
    "1111101011000000",
    "1111101000000001",
    "1111101001010101",
    "1111110010101010",
    "1111111010111010",
    "1111100010000110",
    "1111001000011010",
    "1110110011011000",
    "1110100111011111",
    "1110100110010011",
    "1110101101101000",
    "1110111001011000",
    "1111000101111011",
    "1111010000111101",
    "1111011001011000",
    "1111011110000111",
    "1111011101111010",
    "1111011000010001",
    "1111001101110101",
    "1111000000011001",
    "1110110010111101",
    "1110101000010110",
    "1110100010000000",
    "1110011111111011",
    "1110100000011110",
    "1110100001000101",
    "1110011111101110",
    "1110011011101111",
    "1110010110001000",
    "1110010000111000",
    "1110001101110010",
    "1110001110010110",
    "1110010011010111",
    "1110011101001100",
    "1110101100000001",
    "1111000000000111",
    "1111011001001100",
    "1111110101100101",
    "1111101110011110",
    "1111011000010101",
    "1111001101000100",
    "1111001111111000",
    "1111100000011010",
    "1111111010100010",
    "1111101000010001",
    "1111001111000111",
    "1110111111001101",
    "1110111010100010",
    "1111000000110101",
    "1111010001001111",
    "1111101010001011",
    "1111110110100100",
    "1111010100010011",
    "1110110011011101",
    "1110011000101101",
    "1110001000000110",
    "1110000011111011",
    "1110001011001010",
    "1110011001110101",
    "1110101010101000",
    "1110111000101111",
    "1111000001000101",
    "1111000100010101",
    "1111000111010110",
    "1111001111111000",
    "1111100001000011",
    "1111111001011100",
    "1111101100010001",
    "1111010110100111",
    "1111001011001010",
    "1111001100100110",
    "1111011001011000",
    "1111101111101000",
    "1111110001011101",
    "1111001011110101",
    "1110100010100100",
    "1101111010110111",
    "1101011011011000",
    "1101001001001001",
    "1101000111001001",
    "1101010100011100",
    "1101101011011001",
    "1110000101010010",
    "1110011110010001",
    "1110110110111110",
    "1111010001111000",
    "1111110000001110",
    "1111101111010010",
    "1111010000111001",
    "1110111010110000",
    "1110110010100001",
    "1110111010000010",
    "1111001101010010",
    "1111100100100000",
    "1111110111100011",
    "1111111110101110",
    "1111111110010101",
    "1111111100011011",
    "1111110110001110",
    "1111110010110011",
    "1111110011011011",
    "1111111000101110",
    "1111111011110010",
    "1111101001111010",
    "1111010010111011",
    "1110111001111101",
    "1110100011100111",
    "1110010100010111",
    "1110001111110110",
    "1110010111001000",
    "1110100110011011",
    "1110110111110010",
    "1111000110101010",
    "1111010001100110",
    "1111011001111111",
    "1111100001111000",
    "1111101010000110",
    "1111110010000100",
    "1111110111010010",
    "1111110101110100",
    "1111101010111010",
    "1111010111010011",
    "1110111110100100",
    "1110100110000001",
    "1110010010111110",
    "1110001000100101",
    "1110000111100010",
    "1110001111010100",
    "1110011111010111",
    "1110110111001011",
    "1111010101100111",
    "1111111000000011",
    "1111100101000101",
    "1111000110010011",
    "1110101111111000",
    "1110100100001011",
    "1110100010100111",
    "1110100111011111",
    "1110101110010010",
    "1110110011111000",
    "1110110111011011",
    "1110111011111101",
    "1111000110111001",
    "1111011100100000",
    "1111111101100100",
    "1111011010000010",
    "1110110010001101",
    "1110010011000101",
    "1110000010101110",
    "1110000010110011",
    "1110010000100111",
    "1110101000001011",
    "1111000101100010",
    "1111100101011011",
    "1111111010110110",
    "1111011110010100",
    "1111000111111111",
    "1110111010011001",
    "1110110111011010",
    "1110111111100011",
    "1111010001010010",
    "1111101001101001",
    "1111111010110100",
    "1111011111011110",
    "1111000110111011",
    "1110110011000000",
    "1110100100101110",
    "1110011100010011",
    "1110011001101011",
    "1110011100010001",
    "1110100011100010",
    "1110110000010100",
    "1111000011110001",
    "1111011110000111",
    "1111111110000101",
    "1111011111011111",
    "1110111111001100",
    "1110100101101010",
    "1110010110110010",
    "1110010011110011",
    "1110011010110100",
    "1110101000011010",
    "1110111000111100",
    "1111001001101010",
    "1111011010000001",
    "1111101100101010",
    "1111111011000000",
    "1111011100000001",
    "1110111001000100",
    "1110011000101000",
    "1110000010010100",
    "1101111100001010",
    "1110001000101000",
    "1110100100010111",
    "1111000111011011",
    "1111101001110101",
    "1111111000101100",
    "1111011111111010",
    "1111001001010001",
    "1110110011011100",
    "1110011111001101",
    "1110001111101001",
    "1110001001101101",
    "1110010010100110",
    "1110101100001010",
    "1111010011010011",
    "1111111111010011",
    "1111010101001000",
    "1110110110001001",
    "1110100110010010",
    "1110100101001001",
    "1110101110111010",
    "1110111101110111",
    "1111001100110011",
    "1111011001010000",
    "1111100101011011",
    "1111110101110111",
    "1111110010101001",
    "1111010100100111",
    "1110110100011101",
    "1110011000100111",
    "1110000110100101",
    "1110000010010101",
    "1110001011101011",
    "1110011101111101",
    "1110110011001000",
    "1111000101101100",
    "1111010011000101",
    "1111011101010110",
    "1111101000011110",
    "1111111000000010",
    "1111110010100100",
    "1111011010001011",
    "1111000011111100",
    "1110110101010011",
    "1110110010010100",
    "1110111011001110",
    "1111001100000010",
    "1111011110111010",
    "1111101110100100",
    "1111111000000001",
    "1111111011000010",
    "1111111000111011",
    "1111110100010010",
    "1111110000111111",
    "1111110010101001",
    "1111111010111110",
    "1111110110101110",
    "1111100101101010",
    "1111010110010101",
    "1111001101001111",
    "1111001110000100",
    "1111011010100000",
    "1111110001011001",
    "1111110001000001",
    "1111010010010100",
    "1110110111110010",
    "1110100101010101",
    "1110011100100011",
    "1110011100100101",
    "1110100010101100",
    "1110101100000010",
    "1110110110001110",
    "1111000000000101",
    "1111001001001110",
    "1111010001011001",
    "1111011000100101",
    "1111011111111010",
    "1111101001010110",
    "1111110110101000",
    "1111110111111101",
    "1111100100010101",
    "1111010001101001",
    "1111000011001000",
    "1110111011100000",
    "1110111011110011",
    "1111000010100111",
    "1111001100101010",
    "1111010101111001",
    "1111011010101010",
    "1111011000100111",
    "1111001110101110",
    "1110111101111111",
    "1110101001011000",
    "1110010100110111",
    "1110000100010101",
    "1101111010001110",
    "1101110111010000",
    "1101111010001001",
    "1110000000011111",
    "1110000111101000",
    "1110001101101101",
    "1110010010001111",
    "1110010110000110",
    "1110011011000001",
    "1110100100010010",
    "1110110110000011",
    "1111010010001010",
    "1111110110111010",
    "1111100000101011",
    "1110111011101101",
    "1110100000011110",
    "1110010010111110",
    "1110010011110001",
    "1110011110110110",
    "1110101110011110",
    "1110111101101000",
    "1111001001100000",
    "1111010010000011",
    "1111011001011011",
    "1111100011010011",
    "1111110011101001",
    "1111110100100110",
    "1111011000100000",
    "1110111101101011",
    "1110101010010100",
    "1110100011000000",
    "1110101001001100",
    "1110111010101101",
    "1111010010101001",
    "1111101011011011",
    "1111111111101000",
    "1111110001100101",
    "1111101011001111",
    "1111101011110000",
    "1111110001001011",
    "1111111001001001",
    "1111111110001001",
    "1111110101111000",
    "1111101110100000",
    "1111101000000110",
    "1111100010110001",
    "1111011111000111",
    "1111011110001101",
    "1111100001010100",
    "1111101001100000",
    "1111110111100101",
    "1111110100011001",
    "1111011100000100",
    "1111000010101111",
    "1110101100110000",
    "1110011101111000",
    "1110010111111100",
    "1110011010011000",
    "1110100010111001",
    "1110101110010111",
    "1110111010111111",
    "1111001010100011",
    "1111100000101110",
    "1111111111101110",
    "1111011001100000",
    "1110110000001010",
    "1110001011011110",
    "1101110010000101",
    "1101101000010011",
    "1101101101011100",
    "1101111100000010",
    "1110001101100001",
    "1110011100010111",
    "1110100110110010",
    "1110110000011100",
    "1110111111000111",
    "1111010111001110",
    "1111111000111100",
    "1111100001001111",
    "1110111111100011",
    "1110101000111111",
    "1110100001010100",
    "1110100110100000",
    "1110110001111101",
    "1110111100010001",
    "1111000000100111",
    "1110111110010100",
    "1110111000001001",
    "1110110001100001",
    "1110101101000111",
    "1110101100010100",
    "1110101110010111",
    "1110110010111001",
    "1110111011111100",
    "1111001011101010",
    "1111100011000110",
    "1111111111001001",
    "1111011111111111",
    "1111000101011010",
    "1110110100110011",
    "1110110000100011",
    "1110110110000110",
    "1110111111100011",
    "1111000110110110",
    "1111000111101101",
    "1111000001101011",
    "1110110111001001",
    "1110101011101111",
    "1110100011010000",
    "1110100000001111",
    "1110100010100100",
    "1110101000011000",
    "1110101110110101",
    "1110110011010101",
    "1110110100111001",
    "1110110100000110",
    "1110110010101100",
    "1110110010101100",
    "1110110101011101",
    "1110111011100011",
    "1111000110011000",
    "1111011000010110",
    "1111110011000010",
    "1111101010011011",
    "1111000100000011",
    "1110011111111111",
    "1110000100011010",
    "1101110110000011",
    "1101110110010011",
    "1110000010000110",
    "1110010011110011",
    "1110100101101110",
    "1110110100000000",
    "1110111101110111",
    "1111000100111011",
    "1111001011011110",
    "1111010011011100",
    "1111011100110011",
    "1111100110001011",
    "1111101111000011",
    "1111111000010010",
    "1111111100110100",
    "1111101111011011",
    "1111100000010010",
    "1111010010000000",
    "1111000111111001",
    "1111000100011111",
    "1111001000001001",
    "1111010000100110",
    "1111011010100101",
    "1111100011001010",
    "1111101000111010",
    "1111101100110111",
    "1111110001011010",
    "1111111000111101",
    "1111111011001000",
    "1111101011110100",
    "1111011011111010",
    "1111001110110000",
    "1111000110110111",
    "1111000100110100",
    "1111000110110010",
    "1111001001011101",
    "1111001001110000",
    "1111000110000001",
    "1110111110101110",
    "1110110101101010",
    "1110101101010100",
    "1110101000001011",
    "1110100111111111",
    "1110101101101011",
    "1110111001000110",
    "1111001001001100",
    "1111011100100110",
    "1111110001011111",
    "1111111010000011",
    "1111100111111010",
    "1111011001001011",
    "1111001101111101",
    "1111000101110110",
    "1111000000000010",
    "1110111011110011",
    "1110111001001110",
    "1110111000111100",
    "1110111011101011",
    "1111000001100110",
    "1111001001110000",
    "1111010011100010",
    "1111100000001100",
    "1111110001101001",
    "1111110111010101",
    "1111011100011011",
    "1111000001111110",
    "1110101101101011",
    "1110100100101110",
    "1110101010100000",
    "1110111110101000",
    "1111011100110011",
    "1111111110101100",
    "1111100010010100",
    "1111001011001001",
    "1110111101110101",
    "1110111010000001",
    "1110111101001110",
    "1111000100000000",
    "1111001011110111",
    "1111010011010111",
    "1111011010001110",
    "1111100000111000",
    "1111100111010111",
    "1111101100111010",
    "1111110000100001",
    "1111110001110001",
    "1111110001011000",
    "1111110001001001",
    "1111110011010001",
    "1111111001110001",
    "1111111010001100",
    "1111101001010101",
    "1111010110001110",
    "1111000100101100",
    "1110111000001001",
    "1110110010010101",
    "1110110010101011",
    "1110110111111100",
    "1111000010011111",
    "1111010010111110",
    "1111101000110001",
    "1111111110111110",
    "1111101001010110",
    "1111011011110011",
    "1111011010000111",
    "1111100101001101",
    "1111111001010011",
    "1111110000110010",
    "1111100000001111",
    "1111011001111101",
    "1111011101110111",
    "1111100101101001",
    "1111101001010011",
    "1111100011000011",
    "1111010001100110",
    "1110111001100111",
    "1110100011000001",
    "1110010101011000",
    "1110010101010101",
    "1110100001111001",
    "1110110101001110",
    "1111001001011001",
    "1111011100011001",
    "1111110000010011",
    "1111110111111111",
    "1111011100001100",
    "1110111111010001",
    "1110100110101100",
    "1110011000110111",
    "1110011010001100",
    "1110101010001001",
    "1111000011010011",
    "1111011101110111",
    "1111110011011001",
    "1111111101001011",
    "1111110000001001",
    "1111100000111011",
    "1111001101010010",
    "1110110110110110",
    "1110100010010010",
    "1110010100101100",
    "1110010001001101",
    "1110010111000001",
    "1110100001111001",
    "1110101101000000",
    "1110110101001011",
    "1110111010011000",
    "1110111110111101",
    "1111000101001101",
    "1111001101101110",
    "1111010111011000",
    "1111011111101100",
    "1111100100010101",
    "1111100100010010",
    "1111100000110110",
    "1111011101101001",
    "1111011110100001",
    "1111100101001110",
    "1111110000010010",
    "1111111100000111",
    "1111111010010011",
    "1111110100000111",
    "1111101111111001",
    "1111101010101011",
    "1111100001100010",
    "1111010011011111",
    "1111000010001011",
    "1110110001100111",
    "1110100110001001",
    "1110100010100100",
    "1110100111001001",
    "1110110010000010",
    "1111000001100110",
    "1111010101010010",
    "1111101100110100",
    "1111111000100011",
    "1111011101010001",
    "1111000100111001",
    "1110110011010010",
    "1110101011100110",
    "1110101110100110",
    "1110111001100011",
    "1111000111101000",
    "1111010100010011",
    "1111011101111010",
    "1111100110011110",
    "1111110001101011",
    "1111111101101110",
    "1111100111100101",
    "1111001110101011",
    "1110110111100010",
    "1110100111000001",
    "1110100000111101",
    "1110100111001001",
    "1110111000111110",
    "1111010011100100",
    "1111110010110100",
    "1111101101111011",
    "1111010011011010",
    "1111000001100001",
    "1110111010100000",
    "1110111101111000",
    "1111001000101000",
    "1111010111001000",
    "1111100111101011",
    "1111111011001100",
    "1111101100111101",
    "1111010000101110",
    "1110110010011100",
    "1110010110011010",
    "1110000001110110",
    "1101111001011011",
    "1101111110110011",
    "1110001111010010",
    "1110100101100100",
    "1110111011100101",
    "1111001100100101",
    "1111010110101000",
    "1111011010010110",
    "1111011001110111",
    "1111011001111010",
    "1111011111111111",
    "1111101111001000",
    "1111111001000101",
    "1111011101001010",
    "1111000011110011",
    "1110110011001000",
    "1110101111010110",
    "1110111001010001",
    "1111001101011011",
    "1111100101100111",
    "1111111011110000",
    "1111110010100001",
    "1111100010100100",
    "1111010000110000",
    "1110111011010001",
    "1110100011011000",
    "1110001101101101",
    "1101111111111101",
    "1101111110110000",
    "1110001011010110",
    "1110100010001011",
    "1110111110011011",
    "1111011100101110",
    "1111111011001011",
    "1111100110011110",
    "1111001001010001",
    "1110101111111011",
    "1110011101010111",
    "1110010100011000",
    "1110010110010000",
    "1110100000111001",
    "1110110000011100",
    "1111000000101100",
    "1111001110000010",
    "1111010110111001",
    "1111011100010100",
    "1111100001101001",
    "1111101010100111",
    "1111111000011011",
    "1111110111010010",
    "1111101000110101",
    "1111100000100011",
    "1111100001011110",
    "1111101011101111",
    "1111111100010000",
    "1111110001111010",
    "1111100011110100",
    "1111011100111100",
    "1111011111000100",
    "1111101010110010",
    "1111111111010101",
    "1111100101101010",
    "1111001000001011",
    "1110101100110000",
    "1110010111011011",
    "1110001010100110",
    "1110000110101111",
    "1110001001111010",
    "1110010000101011",
    "1110010111000100",
    "1110011010101010",
    "1110011100111101",
    "1110100011100001",
    "1110110011111011",
    "1111010000010101",
    "1111110101111001",
    "1111100010011010",
    "1111000000100110",
    "1110101010111010",
    "1110100011100111",
    "1110100111100011",
    "1110110000100100",
    "1110111000101111",
    "1110111100100101",
    "1110111100001110",
    "1110111001110010",
    "1110110111110111",
    "1110111000011011",
    "1110111100000100",
    "1111000001100100",
    "1111000110111110",
    "1111001010101111",
    "1111001100100110",
    "1111001101010110",
    "1111001101101101",
    "1111001101101011",
    "1111001100011110",
    "1111001001100000",
    "1111000101010010",
    "1111000001100010",
    "1111000000110001",
    "1111000101011111",
    "1111010001011110",
    "1111100101001011",
    "1111111111011100",
    "1111100010101001",
    "1111000100110100",
    "1110101010011011",
    "1110010110001001",
    "1110001001101010",
    "1110000101100111",
    "1110001001011011",
    "1110010011010101",
    "1110100000101110",
    "1110101110110011",
    "1110111010101010",
    "1111000010100100",
    "1111001000110100",
    "1111010010100010",
    "1111100011110100",
    "1111111101100101",
    "1111100011110110",
    "1111000111011000",
    "1110110011110011",
    "1110101101111011",
    "1110110101111011",
    "1111000110101111",
    "1111011001111001",
    "1111101001101001",
    "1111110100000010",
    "1111111100010001",
    "1111111000110000",
    "1111100111110101",
    "1111010000111101",
    "1110111000101000",
    "1110100101010011",
    "1110011100001100",
    "1110011111101001",
    "1110101101100011",
    "1111000000100100",
    "1111010011001111",
    "1111100010000110",
    "1111101100111111",
    "1111110101100101",
    "1111111101011010",
    "1111111010101010",
    "1111110010110011",
    "1111101100010111",
    "1111101000110010",
    "1111101001000111",
    "1111101101101010",
    "1111110101100110",
    "1111111111101101",
    "1111110100010101",
    "1111100110000000",
    "1111010100011010",
    "1110111111110110",
    "1110101010011001",
    "1110010111011000",
    "1110001010010100",
    "1110000101110110",
    "1110001010100011",
    "1110010110111011",
    "1110100111111100",
    "1110111010010001",
    "1111001011000111",
    "1111011000101101",
    "1111100001111001",
    "1111100110010000",
    "1111100101110001",
    "1111100001001010",
    "1111011001110111",
    "1111010001111000",
    "1111001011011110",
    "1111001001000010",
    "1111001100010111",
    "1111010101110110",
    "1111100011111000",
    "1111110011100100",
    "1111111101111000",
    "1111110010001111",
    "1111101001010110",
    "1111100001011110",
    "1111011000010101",
    "1111001100100110",
    "1110111110101001",
    "1110110000011111",
    "1110100100110110",
    "1110011101110010",
    "1110011011110010",
    "1110011101100100",
    "1110100000110001",
    "1110100011010011",
    "1110100100010111",
    "1110100100011101",
    "1110100110101000",
    "1110101111100001",
    "1111000010010010",
    "1111011110011001",
    "1111111111011100",
    "1111100001100001",
    "1111001011001001",
    "1111000010000011",
    "1111000111111001",
    "1111011010010100",
    "1111110100100000",
    "1111101111000010",
    "1111010101011000",
    "1111000001110000",
    "1110110101110001",
    "1110110010000101",
    "1110110101110110",
    "1110111111011111",
    "1111001101001010",
    "1111011100111010",
    "1111101101000111",
    "1111111100011101",
    "1111110110000001",
    "1111101010110001",
    "1111100001100110",
    "1111011001111010",
    "1111010011011010",
    "1111001110011011",
    "1111001011101011",
    "1111001011110010",
    "1111001110101011",
    "1111010011101110",
    "1111011001111111",
    "1111100000100100",
    "1111100110111011",
    "1111101100100100",
    "1111110001101001",
    "1111111000001010",
    "1111111100110000",
    "1111101011100111",
    "1111010101100111",
    "1110111110100011",
    "1110101011011011",
    "1110100000011100",
    "1110011111110110",
    "1110101000101000",
    "1110110110011101",
    "1111000100010010",
    "1111001110001111",
    "1111010010110110",
    "1111010010111000",
    "1111001111111011",
    "1111001011010100",
    "1111000101100101",
    "1110111110011110",
    "1110110101100100",
    "1110101011000110",
    "1110100000000111",
    "1110010110100101",
    "1110010000100111",
    "1110001111010010",
    "1110010001110100",
    "1110010110101100",
    "1110011110110001",
    "1110101101001010",
    "1111000100010010",
    "1111100100001101",
    "1111110110010111",
    "1111010001010100",
    "1110110010101100",
    "1110011111011010",
    "1110011000111010",
    "1110011100001001",
    "1110100100001000",
    "1110101100000100",
    "1110110001000111",
    "1110110011100010",
    "1110110101000110",
    "1110111000001100",
    "1110111111110101",
    "1111001101111010",
    "1111100010001000",
    "1111111010001111",
    "1111101101110001",
    "1111011001111111",
    "1111001100111100",
    "1111000111011000",
    "1111001000001011",
    "1111001100011001",
    "1111010000100001",
    "1111010001101001",
    "1111001110101110",
    "1111001001011110",
    "1111000101001101",
    "1111000101100010",
    "1111001100111100",
    "1111011011010110",
    "1111101110001110",
    "1111111110010100",
    "1111101110101000",
    "1111100101100101",
    "1111100011111001",
    "1111101000001001",
    "1111101111111011",
    "1111111000111011",
    "1111111110011101",
    "1111110111011011",
    "1111110010011101",
    "1111101111100000",
    "1111101110011100",
    "1111101111000101",
    "1111110001000110",
    "1111110100000010",
    "1111110111000001",
    "1111111001000010",
    "1111111001011110",
    "1111111000011011",
    "1111110110110001",
    "1111110101101001",
    "1111110110000011",
    "1111111000101101",
    "1111111101110000",
    "1111111011001111",
    "1111110011001100",
    "1111101010111011",
    "1111100011001101",
    "1111011100111100",
    "1111011001011000",
    "1111011001111111",
    "1111011111100011",
    "1111101001110010",
    "1111110110111111",
    "1111111011010111",
    "1111110000000100",
    "1111101001000101",
    "1111100111010001",
    "1111101010001000",
    "1111110000011110",
    "1111111001000000",
    "1111111101001110",
    "1111110010101100",
    "1111100111111011",
    "1111011101101011",
    "1111010101000110",
    "1111001111001100",
    "1111001100011100",
    "1111001100101010",
    "1111001110110011",
    "1111010001001100",
    "1111010010010101",
    "1111010001100110",
    "1111001111101001",
    "1111001110010100",
    "1111001111110110",
    "1111010110100000",
    "1111100011110100",
    "1111110111101010",
    "1111101111111001",
    "1111010110100100",
    "1111000000101001",
    "1110110001110110",
    "1110101100001010",
    "1110101111011010",
    "1110111001001011",
    "1111000101110110",
    "1111010001110001",
    "1111011010010011",
    "1111011110011011",
    "1111011110011001",
    "1111011011011000",
    "1111010110110010",
    "1111010010001011",
    "1111001110111101",
    "1111001110001100",
    "1111010000110001",
    "1111010111000110",
    "1111100000101100",
    "1111101100011101",
    "1111111000100010",
    "1111111101000111",
    "1111110110000101",
    "1111110011001000",
    "1111110100000000",
    "1111110111101101",
    "1111111101000100",
    "1111111100101100",
    "1111110101101001",
    "1111101101010001",
    "1111100011010011",
    "1111011000010001",
    "1111001101001100",
    "1111000011011101",
    "1110111100001010",
    "1110110111101101",
    "1110110101100101",
    "1110110100101110",
    "1110110100000101",
    "1110110011011101",
    "1110110011100001",
    "1110110101100101",
    "1110111101001010",
    "1111001110011011",
    "1111101011000010",
    "1111101110100010",
    "1111000011101010",
    "1110011011100011",
    "1101111100110011",
    "1101101100000101",
    "1101101010000001",
    "1101110010100110",
    "1110000000000111",
    "1110001101000101",
    "1110010101100111",
    "1110011000100010",
    "1110010110010000",
    "1110010000010101",
    "1110001001001110",
    "1110000010101011",
    "1101111110000100",
    "1101111110010001",
    "1110000110110100",
    "1110011010000001",
    "1110110111011101",
    "1111011011010110",
    "1111111111001111",
    "1111100011011000",
    "1111010001101011",
    "1111001101001010",
    "1111010100001011",
    "1111100011101111",
    "1111111000010110",
    "1111110001011011",
    "1111011100100011",
    "1111001011110011",
    "1111000001100001",
    "1110111111000010",
    "1111000100111100",
    "1111010010110011",
    "1111100110101001",
    "1111111101101001",
    "1111101011101010",
    "1111011001001110",
    "1111001110001111",
    "1111001100000101",
    "1111010001101110",
    "1111011100001111",
    "1111101000010100",
    "1111110011100100",
    "1111111100111111",
    "1111111010011010",
    "1111110000010001",
    "1111100001111110",
    "1111001110000101",
    "1110110101010011",
    "1110011010111010",
    "1110000011101110",
    "1101110100011101",
    "1101110000000111",
    "1101110110100010",
    "1110000101010011",
    "1110011000110111",
    "1110101101110101",
    "1111000011110110",
    "1111011101100100",
    "1111111101001000",
    "1111011101110011",
    "1110110111001101",
    "1110010101110001",
    "1101111111111101",
    "1101111010001110",
    "1110000100111110",
    "1110011011001111",
    "1110110101011101",
    "1111001100101110",
    "1111011101011110",
    "1111101001001011",
    "1111110011110111",
    "1111111111000001",
    "1111101110001100",
    "1111011011101010",
    "1111001011110000",
    "1111000010011111",
    "1111000010010010",
    "1111001010110010",
    "1111011000111100",
    "1111101000110111",
    "1111110111100010",
    "1111111100010111",
    "1111110011010011",
    "1111101101110000",
    "1111101100110100",
    "1111110001100100",
    "1111111100110001",
    "1111110001111000",
    "1111011100100000",
    "1111000110100100",
    "1110110100001011",
    "1110101000111110",
    "1110100110101100",
    "1110101101000111",
    "1110111011010110",
    "1111010000110001",
    "1111101100111011",
    "1111110001011111",
    "1111001101010110",
    "1110101010100110",
    "1110001101110010",
    "1101111010101000",
    "1101110011000101",
    "1101110110001110",
    "1110000000110000",
    "1110001110001010",
    "1110011011000110",
    "1110100111110111",
    "1110110111110100",
    "1111001110100001",
    "1111101101001011",
    "1111101110101110",
    "1111001010111111",
    "1110101110011110",
    "1110011110100110",
    "1110011100111111",
    "1110100110001110",
    "1110110100000001",
    "1111000001101110",
    "1111001111010001",
    "1111011111101110",
    "1111110101110110",
    "1111101110010001",
    "1111010000000111",
    "1110110101100101",
    "1110100110000001",
    "1110100111110100",
    "1110111100101101",
    "1111100000101100",
    "1111110100010001",
    "1111001011111100",
    "1110101101111000",
    "1110011101111010",
    "1110011100010011",
    "1110100101110100",
    "1110110101011011",
    "1111000111110010",
    "1111011100010110",
    "1111110100010010",
    "1111101111101110",
    "1111010001100001",
    "1110110100110111",
    "1110011101111010",
    "1110001111101001",
    "1110001011001100",
    "1110001111001100",
    "1110011000111001",
    "1110100101000000",
    "1110110000111011",
    "1110111011110011",
    "1111000110001000",
    "1111010000011100",
    "1111011010110100",
    "1111100100011010",
    "1111101100000000",
    "1111110010011111",
    "1111111011000100",
    "1111110111101011",
    "1111100101100000",
    "1111010001000000",
    "1110111111010111",
    "1110110101110001",
    "1110110111110001",
    "1111000101001000",
    "1111011000101111",
    "1111101011111100",
    "1111111001010110",
    "1111111110101000",
    "1111111100110100",
    "1111110111100011",
    "1111110101000101",
    "1111111100000000",
    "1111110000110101",
    "1111010011100100",
    "1110110010011010",
    "1110010101001011",
    "1110000010001111",
    "1101111100101110",
    "1110000011100010",
    "1110010010001010",
    "1110100011100110",
    "1110110011110100",
    "1111000000011010",
    "1111001001001001",
    "1111001110101011",
    "1111010010001101",
    "1111010100101111",
    "1111010110011000",
    "1111010110110010",
    "1111010101100101",
    "1111010010100100",
    "1111001110010100",
    "1111001010001100",
    "1111001000001100",
    "1111001010111100",
    "1111010101000000",
    "1111100111110111",
    "1111111100111001",
    "1111011100100011",
    "1110111100100110",
    "1110100011000001",
    "1110010100001000",
    "1110010000110110",
    "1110010110001001",
    "1110011111001100",
    "1110100111010011",
    "1110101011100001",
    "1110101011100000",
    "1110101000110101",
    "1110100111011000",
    "1110101100110010",
    "1110111101010110",
    "1111011001101111",
    "1111111110010011",
    "1111011100001010",
    "1110111101110011",
    "1110101100111101",
    "1110101101000010",
    "1110111101000000",
    "1111011000100010",
    "1111111010000000",
    "1111100100000001",
    "1111000101100101",
    "1110101100110111",
    "1110011011001111",
    "1110010001001101",
    "1110001111001100",
    "1110010110001001",
    "1110100110110100",
    "1111000000011001",
    "1111100000001100",
    "1111111110001011",
    "1111011111100100",
    "1111000111110111",
    "1110111000111010",
    "1110110010100010",
    "1110110010111101",
    "1110110111101101",
    "1110111110010001",
    "1111000100111001",
    "1111001100001100",
    "1111010110110001",
    "1111100111010000",
    "1111111110011110",
    "1111100101111100",
    "1111001010111111",
    "1110110110000110",
    "1110101011110000",
    "1110101101100000",
    "1110111010101101",
    "1111010010101100",
    "1111110100000000",
    "1111100100000110",
    "1110111010000010",
    "1110010011111110",
    "1101111000001110",
    "1101101011011101",
    "1101101111110011",
    "1110000011000101",
    "1110011111111101",
    "1111000010011010",
    "1111101000101001",
    "1111101110011110",
    "1111000100110011",
    "1110011101101001",
    "1101111101001110",
    "1101100111001110",
    "1101011111000101",
    "1101100101010010",
    "1101110101110010",
    "1110001010100011",
    "1110011101100001",
    "1110101010110101",
    "1110110010100010",
    "1110110110110111",
    "1110111010101101",
    "1111000000011111",
    "1111001000011010",
    "1111010010101110",
    "1111100001110001",
    "1111110111000100",
    "1111101101101101",
    "1111001111001101",
    "1110110010101110",
    "1110011101110101",
    "1110010101001000",
    "1110011010011001",
    "1110101010001011",
    "1110111101110000",
    "1111001110101001",
    "1111011000000001",
    "1111011000100000",
    "1111010001111011",
    "1111000111100000",
    "1110111110110011",
    "1110111101110101",
    "1111000111110101",
    "1111011100101000",
    "1111111000010100",
    "1111101011011100",
    "1111010100101110",
    "1111000111110001",
    "1111000110001011",
    "1111001101111011",
    "1111011010110000",
    "1111100111110010",
    "1111110000110110",
    "1111110100010101",
    "1111110010111101",
    "1111101110100001",
    "1111101001100100",
    "1111100101111100",
    "1111100100001000",
    "1111100011101110",
    "1111100011101110",
    "1111100011010000",
    "1111100010101110",
    "1111100011100110",
    "1111100111101101",
    "1111110000011000",
    "1111111110000010",
    "1111101111111001",
    "1111011011011001",
    "1111000111011010",
    "1110110110101000",
    "1110101010111100",
    "1110100100111100",
    "1110100100100100",
    "1110101001101011",
    "1110110100110111",
    "1111000110100111",
    "1111011110100011",
    "1111111010111111",
    "1111100111000000",
    "1111001010111000",
    "1110110011101010",
    "1110100011011000",
    "1110011010011001",
    "1110010111110001",
    "1110011010101101",
    "1110100011101110",
    "1110110011111110",
    "1111001011110011",
    "1111101001100111",
    "1111110110010100",
    "1111011000111110",
    "1111000011000011",
    "1110110111111001",
    "1110111000000100",
    "1111000001011111",
    "1111010000101100",
    "1111100010010010",
    "1111110011111010",
    "1111111011110000",
    "1111101101110000",
    "1111100011010101",
    "1111011101111010",
    "1111011111000000",
    "1111100111110100",
    "1111111000010111",
    "1111110000101101",
    "1111010110010010",
    "1110111011111000",
    "1110100100101010",
    "1110010010110001",
    "1110000111010110",
    "1110000010111110",
    "1110000101110111",
    "1110010000001000",
    "1110100001101001",
    "1110111001101011",
    "1111010110101100",
    "1111110110010111",
    "1111101001111001",
    "1111001100101000",
    "1110110011011111",
    "1110011111010001",
    "1110010000011110",
    "1110000111100000",
    "1110000100111110",
    "1110001001001001",
    "1110010011111001",
    "1110100101100010",
    "1110111111001100",
    "1111100000111000",
    "1111110111100010",
    "1111001110010111",
    "1110101001000110",
    "1110001100110111",
    "1101111101001010",
    "1101111010111111",
    "1110000100000001",
    "1110010011100100",
    "1110100101001011",
    "1110110111100011",
    "1111001100011100",
    "1111100101110010",
    "1111111100011111",
    "1111011101010111",
    "1111000001111101",
    "1110101111111000",
    "1110101011111010",
    "1110110111110111",
    "1111010001100001",
    "1111110011010111",
    "1111101001110100",
    "1111001100110101",
    "1110111001111010",
    "1110110011001111",
    "1110111000110010",
    "1111001000011101",
    "1111011110110101",
    "1111111000000111",
    "1111101111010001",
    "1111011010001001",
    "1111001010011110",
    "1111000001111001",
    "1111000001001000",
    "1111000111011010",
    "1111010010101011",
    "1111100000011111",
    "1111101110100001",
    "1111111010101001",
    "1111111100111010",
    "1111111001001000",
    "1111111001110000",
    "1111111101100101",
    "1111111101010100",
    "1111111001001100",
    "1111111000001011",
    "1111111100000111",
    "1111111010000011",
    "1111101010111011",
    "1111011000011101",
    "1111000101101111",
    "1110110110000011",
    "1110101100000111",
    "1110101001001011",
    "1110101100101000",
    "1110110100010000",
    "1110111101001001",
    "1111000100101110",
    "1111001001100111",
    "1111001011101010",
    "1111001011101101",
    "1111001010111000",
    "1111001010011011",
    "1111001011001111",
    "1111001110000101",
    "1111010100110100",
    "1111100010010000",
    "1111110111111101",
    "1111101010101100",
    "1111001001010101",
    "1110101001111010",
    "1110010010011101",
    "1110000111100010",
    "1110001010001001",
    "1110010111000001",
    "1110101000110010",
    "1110111010111010",
    "1111001010101111",
    "1111011000000001",
    "1111100011100001",
    "1111101101011000",
    "1111110101001011",
    "1111111001100110",
    "1111111001010101",
    "1111110100101111",
    "1111101110000011",
    "1111101000101111",
    "1111101000001110",
    "1111101110011001",
    "1111111010100101",
    "1111110110010100",
    "1111101000110011",
    "1111100000100001",
    "1111011111000101",
    "1111100011101001",
    "1111101011100100",
    "1111110011010010",
    "1111110111101011",
    "1111110111010000",
    "1111110011001100",
    "1111101111000010",
    "1111101110110001",
    "1111110101001110",
    "1111111100111110",
    "1111101001101001",
    "1111010100000110",
    "1111000000001101",
    "1110110000110101",
    "1110100110110010",
    "1110100001010100",
    "1110011111001010",
    "1110011111010001",
    "1110100001000111",
    "1110100100100100",
    "1110101001011101",
    "1110101111001111",
    "1110110101000001",
    "1110111001010000",
    "1110111010011101",
    "1110110111101111",
    "1110110001000101",
    "1110100111101100",
    "1110011101101000",
    "1110010101010111",
    "1110010001111000",
    "1110010101101100",
    "1110100001101011",
    "1110110011111110",
    "1111001000000110",
    "1111011000010101",
    "1111011111111101",
    "1111011100111111",
    "1111010001000010",
    "1111000000111101",
    "1110110010110001",
    "1110101100000101",
    "1110110000011111",
    "1111000000110000",
    "1111011010101011",
    "1111111001111100",
    "1111100110110110",
    "1111001100111010",
    "1110111100010001",
    "1110110111000100",
    "1110111101001100",
    "1111001100101011",
    "1111100010010100",
    "1111111010001000",
    "1111101111110011",
    "1111011111000100",
    "1111010110000011",
    "1111010101101111",
    "1111011101100100",
    "1111101011111001",
    "1111111110001000",
    "1111101110101101",
    "1111011101111010",
    "1111010010100001",
    "1111001110101001",
    "1111010010100110",
    "1111011100101010",
    "1111101001100100",
    "1111110101011111",
    "1111111100111101",
    "1111111101101100",
    "1111110110111010",
    "1111101001011000",
    "1111010111010000",
    "1111000011101001",
    "1110110010000011",
    "1110100101011101",
    "1110011111011110",
    "1110100000000000",
    "1110100110001101",
    "1110110001111101",
    "1111000011011111",
    "1111011010001001",
    "1111110011101010",
    "1111110011110011",
    "1111100000110000",
    "1111010110010000",
    "1111010101011000",
    "1111011100001111",
    "1111100110100100",
    "1111101111110011",
    "1111110100110000",
    "1111110100100100",
    "1111110000111000",
    "1111101100111101",
    "1111101101001110",
    "1111110101100101",
    "1111111000110010",
    "1111100000001101",
    "1111000101100000",
    "1110101110110001",
    "1110100001010000",
    "1110011111111111",
    "1110101010111100",
    "1110111111010111",
    "1111011001000111",
    "1111110011011111",
    "1111110101110011",
    "1111100110000000",
    "1111011110111000",
    "1111100001001010",
    "1111101100101111",
    "1111111111010100",
    "1111100101001101",
    "1111001000000110",
    "1110101011111010",
    "1110010100110110",
    "1110000110011000",
    "1110000010001011",
    "1110000111100011",
    "1110010011100110",
    "1110100010111101",
    "1110110011101001",
    "1111000101000110",
    "1111010111011011",
    "1111101010011101",
    "1111111101010000",
    "1111110001110100",
    "1111100100100100",
    "1111011100001001",
    "1111011000001110",
    "1111010110111100",
    "1111010101110110",
    "1111010011010000",
    "1111001111001100",
    "1111001011001100",
    "1111001001100000",
    "1111001011110000",
    "1111010010010000",
    "1111011011101000",
    "1111100101011101",
    "1111101101001101",
    "1111110000111110",
    "1111110000000100",
    "1111101010111100",
    "1111100010101100",
    "1111011000100111",
    "1111001110010111",
    "1111000111000100",
    "1111000111000011",
    "1111010001101100",
    "1111100111110101",
    "1111111001010100",
    "1111010111011101",
    "1110111001010000",
    "1110100100001110",
    "1110011010111101",
    "1110011011111100",
    "1110100011000011",
    "1110101011101000",
    "1110110010010100",
    "1110110110000110",
    "1110110111100101",
    "1110110111111100",
    "1110111000010110",
    "1110111001000110",
    "1110111001110000",
    "1110111010101010",
    "1110111101110011",
    "1111000101110110",
    "1111010100101010",
    "1111101001100101",
    "1111111111011010",
    "1111101100100111",
    "1111100100100010",
    "1111101011011100",
    "1111111110101001",
    "1111011110001100",
    "1110111010010001",
    "1110011010101111",
    "1110000101011111",
    "1101111101001110",
    "1110000001001100",
    "1110001101101000",
    "1110011110101110",
    "1110110011101001",
    "1111001101001110",
    "1111101011111101",
    "1111110001011000",
    "1111001111000000",
    "1110110010011010",
    "1110100000100011",
    "1110011011111100",
    "1110100010110011",
    "1110101111111011",
    "1110111101011001",
    "1111000110100100",
    "1111001001011001",
    "1111000110110010",
    "1111000000110011",
    "1110111010110000",
    "1110111001101000",
    "1111000001111110",
    "1111010101101010",
    "1111110011000000",
    "1111101011011001",
    "1111001100101010",
    "1110110111000100",
    "1110101111000000",
    "1110110101000001",
    "1111000101010000",
    "1111011001001001",
    "1111101001110110",
    "1111110010110101",
    "1111110011001101",
    "1111101110000010",
    "1111101001111100",
    "1111101101101010",
    "1111111011111010",
    "1111101101011101",
    "1111010100100010",
    "1111000000011001",
    "1110110110011111",
    "1110111001000111",
    "1111000110101100",
    "1111011011010011",
    "1111110011001111",
    "1111110100100000",
    "1111011110000100",
    "1111001010110101",
    "1110111100011011",
    "1110110100010011",
    "1110110011110011",
    "1110111011111111",
    "1111001101000000",
    "1111100101100111",
    "1111111100100000",
    "1111011100100011",
    "1110111101101001",
    "1110100010011101",
    "1110001100110010",
    "1101111101111111",
    "1101110110111100",
    "1101111000000100",
    "1110000001011110",
    "1110010011010101",
    "1110101101011100",
    "1111001110001001",
    "1111110010001001",
    "1111101010111000",
    "1111001101100110",
    "1110111001101000",
    "1110110000110001",
    "1110110001111110",
    "1110111001100101",
    "1111000010111110",
    "1111001010100110",
    "1111001111000111",
    "1111010001000111",
    "1111010010000011",
    "1111010011010101",
    "1111010101101010",
    "1111011000110100",
    "1111011011101111",
    "1111011101010001",
    "1111011100101101",
    "1111011001110100",
    "1111010101001000",
    "1111001111011100",
    "1111001001100111",
    "1111000100011100",
    "1111000000100110",
    "1110111110110000",
    "1111000000100110",
    "1111001001000100",
    "1111011010100010",
    "1111110101010000",
    "1111101001000001",
    "1111000100110001",
    "1110100011010010",
    "1110001001011101",
    "1101111010010110",
    "1101110101110110",
    "1101111001010110",
    "1110000001001111",
    "1110001010000100",
    "1110010001101100",
    "1110010111011011",
    "1110011011110010",
    "1110100000010101",
    "1110100110111011",
    "1110110000110110",
    "1110111110101101",
    "1111001111110101",
    "1111100010011100",
    "1111110100000011",
    "1111111101110100",
    "1111110101011010",
    "1111110011110001",
    "1111111000101111",
    "1111111100111101",
    "1111101111001011",
    "1111011111011010",
    "1111001110111010",
    "1110111111000101",
    "1110110001110001",
    "1110101010001011",
    "1110101100011100",
    "1110111011110101",
    "1111011000010011",
    "1111111101111100",
    "1111011010010110",
    "1110111000110010",
    "1110100011111001",
    "1110011110101011",
    "1110100111101100",
    "1110111001110101",
    "1111010000001101",
    "1111101001010101",
    "1111111001110011",
    "1111011000011110",
    "1110110011111110",
    "1110010000100100",
    "1101110100001010",
    "1101100100001101",
    "1101100011101111",
    "1101110000110110",
    "1110000101010101",
    "1110011010001100",
    "1110101001111001",
    "1110110010101100",
    "1110111000011110",
    "1111000010101110",
    "1111010111110001",
    "1111111001101100",
    "1111011011101011",
    "1110110001001010",
    "1110001111111000",
    "1101111110111010",
    "1110000000011010",
    "1110010000010100",
    "1110100111100011",
    "1110111111011100",
    "1111010011010000",
    "1111100001010000",
    "1111101001011101",
    "1111101100110101",
    "1111101110010001",
    "1111110001010011",
    "1111111000100101",
    "1111111010100010",
    "1111101001001111",
    "1111010110110010",
    "1111000111001011",
    "1110111101111111",
    "1110111101001010",
    "1111000011110001",
    "1111001110011110",
    "1111011000100111",
    "1111011110001010",
    "1111011101100001",
    "1111010111101111",
    "1111001111100100",
    "1111001000001110",
    "1111000011100111",
    "1111000001110001",
    "1111000001011001",
    "1111000000111001",
    "1110111111101000",
    "1110111111001010",
    "1111000011011111",
    "1111010000111011",
    "1111101001101001",
    "1111110011110010",
    "1111001100011100",
    "1110100110111111",
    "1110001001111001",
    "1101111001000100",
    "1101110100100101",
    "1101111001001100",
    "1110000010011100",
    "1110001100100001",
    "1110010101100010",
    "1110011101011100",
    "1110100100111011",
    "1110101100101011",
    "1110110100111110",
    "1110111110111111",
    "1111001101010001",
    "1111100001110000",
    "1111111100100100",
    "1111100100001010",
    "1111000100100010",
    "1110101001011001",
    "1110010111011101",
    "1110010001001101",
    "1110010101101010",
    "1110100001111001",
    "1110110011000101",
    "1111000111011011",
    "1111011110000010",
    "1111110101101011",
    "1111110011110001",
    "1111100000111110",
    "1111010100100101",
    "1111010000010100",
    "1111010011101110",
    "1111011100100001",
    "1111100111011010",
    "1111110001001011",
    "1111110111110101",
    "1111111010111110",
    "1111111011001011",
    "1111111001010100",
    "1111110101101010",
    "1111101111111100",
    "1111100111110010",
    "1111011101010001",
    "1111010001000111",
    "1111000100101001",
    "1110111001101010",
    "1110110001101001",
    "1110101101100100",
    "1110101101101001",
    "1110110001101001",
    "1110111001011000",
    "1111000100110001",
    "1111010011100110",
    "1111100101001110",
    "1111111000110001",
    "1111110010111110",
    "1111011111011110",
    "1111001110010110",
    "1111000001000000",
    "1110111000010000",
    "1110110011111110",
    "1110110011100100",
    "1110110110010110",
    "1110111100001110",
    "1111000110000110",
    "1111010110000001",
    "1111101101100111",
    "1111110011010010",
    "1111001111011111",
    "1110101011110010",
    "1110001101101110",
    "1101111001111001",
    "1101110010011001",
    "1101110110000110",
    "1110000001011010",
    "1110001111110110",
    "1110011101011110",
    "1110100111111100",
    "1110101111111011",
    "1110111010000001",
    "1111001011100011",
    "1111100110111110",
    "1111110101011011",
    "1111001111011100",
    "1110101110010001",
    "1110011000011110",
    "1110010010010101",
    "1110011011110111",
    "1110110001010010",
    "1111001101001001",
    "1111101001010000",
    "1111111111110011",
    "1111110010010011",
    "1111110001001101",
    "1111111101001000",
    "1111101100000101",
    "1111001110101110",
    "1110110000100011",
    "1110010111011101",
    "1110000111100111",
    "1110000010101111",
    "1110001000000011",
    "1110010100010111",
    "1110100011011111",
    "1110110001110110",
    "1110111101110101",
    "1111000111110101",
    "1111010000111101",
    "1111011001101111",
    "1111100001111101",
    "1111101000110001",
    "1111101101011100",
    "1111101111110110",
    "1111110000010011",
    "1111101111100111",
    "1111101110110011",
    "1111101110110111",
    "1111110000011001",
    "1111110011110010",
    "1111111001001100",
    "1111111111100000",
    "1111110110111011",
    "1111101110000000",
    "1111100101100101",
    "1111011110011011",
    "1111011001000001",
    "1111010101100111",
    "1111010011111100",
    "1111010011000110",
    "1111010001111101",
    "1111001111101001",
    "1111001100001001",
    "1111001001001001",
    "1111001001100101",
    "1111010000000111",
    "1111011101100011",
    "1111110000001011",
    "1111111011101111",
    "1111101011001010",
    "1111100010011101",
    "1111100011110100",
    "1111101110010011",
    "1111111110101101",
    "1111101110111010",
    "1111011110000111",
    "1111010001001101",
    "1111001001100010",
    "1111000111010001",
    "1111001001110010",
    "1111001111111101",
    "1111011000011010",
    "1111100001011100",
    "1111101001000101",
    "1111101101110000",
    "1111101110100100",
    "1111101011110010",
    "1111100111000111",
    "1111100011001010",
    "1111100010110011",
    "1111101000011000",
    "1111110100111101",
    "1111111000000010",
    "1111100001000000",
    "1111001001100000",
    "1110110101100111",
    "1110101000110010",
    "1110100100111011",
    "1110101001101101",
    "1110110100111011",
    "1111000011000101",
    "1111010000100100",
    "1111011010100011",
    "1111011111101110",
    "1111100000100100",
    "1111011110110011",
    "1111011100100110",
    "1111011100100000",
    "1111100010110001",
    "1111110011011101",
    "1111110000001111",
    "1111001010101101",
    "1110100001110011",
    "1101111100111100",
    "1101100010101111",
    "1101010111011011",
    "1101011010111010",
    "1101101000110100",
    "1101111011011000",
    "1110001101001111",
    "1110011011001100",
    "1110100100101001",
    "1110101010011000",
    "1110101110001001",
    "1110110001100110",
    "1110110110000000",
    "1110111101110101",
    "1111001011111101",
    "1111100001010101",
    "1111111100100000",
    "1111100110100101",
    "1111001101101110",
    "1110111111000111",
    "1110111111111111",
    "1111010001011100",
    "1111101111011110",
    "1111101100110111",
    "1111001011010110",
    "1110110010011101",
    "1110100110111110",
    "1110101011111010",
    "1111000001001100",
    "1111100011001010",
    "1111110100001111",
    "1111001100100001",
    "1110101100101101",
    "1110011001111001",
    "1110010110000110",
    "1110011111111010",
    "1110110010111000",
    "1111001001010101",
    "1111011110001001",
    "1111101101110111",
    "1111111000001100",
    "1111111111000111",
    "1111110011000110",
    "1111100000101011",
    "1111001000011010",
    "1110101110110000",
    "1110011001110000",
    "1110001110100001",
    "1110001111011010",
    "1110011010011101",
    "1110101010011011",
    "1110111010011001",
    "1111000111010101",
    "1111010000101110",
    "1111011000001110",
    "1111011111101001",
    "1111101000001100",
    "1111110001011011",
    "1111111001010100",
    "1111111110101110",
    "1111111100110010",
    "1111110110100110",
    "1111101100011101",
    "1111011101111111",
    "1111001101010110",
    "1110111110010111",
    "1110110101000110",
    "1110110011110001",
    "1110111001001011",
    "1111000001111001",
    "1111001011101101",
    "1111010111010000",
    "1111100111001101",
    "1111111101111111",
    "1111100100101111",
    "1111000100101100",
    "1110100111100000",
    "1110010011011111",
    "1110001100101110",
    "1110010011001010",
    "1110100010111001",
    "1110110110000001",
    "1111000111001001",
    "1111010101011010",
    "1111100100000000",
    "1111110111000111",
    "1111101110111111",
    "1111010000000111",
    "1110110001010010",
    "1110011000100000",
    "1110001010100010",
    "1110001000111001",
    "1110010001100001",
    "1110100000110110",
    "1110110011101110",
    "1111000111111110",
    "1111011100011011",
    "1111101111011000",
    "1111111110100000",
    "1111111000011011",
    "1111110111001011",
    "1111111110000010",
    "1111110100110110",
    "1111100101001011",
    "1111010111010110",
    "1111001111010110",
    "1111001111001010",
    "1111010110010110",
    "1111100010100010",
    "1111110001000010",
    "1111111111111100",
    "1111110001100111",
    "1111100100000000",
    "1111010111100010",
    "1111001100101110",
    "1111000100001110",
    "1110111110010110",
    "1110111010101011",
    "1110111000010101",
    "1110110110001011",
    "1110110011101001",
    "1110110001011001",
    "1110110010000101",
    "1110111001111010",
    "1111001100001001",
    "1111101001010101",
    "1111110001011000",
    "1111001001100111",
    "1110100101101010",
    "1110001010111000",
    "1101111011101011",
    "1101110110111100",
    "1101111001100010",
    "1110000000000000",
    "1110000111101101",
    "1110001111000111",
    "1110010101010011",
    "1110011001101010",
    "1110011100000101",
    "1110011101000000",
    "1110011101011011",
    "1110011110111011",
    "1110100011010111",
    "1110101011111101",
    "1110111000111100",
    "1111001000110100",
    "1111011000101101",
    "1111100101110001",
    "1111101110110011",
    "1111110101001001",
    "1111111011110011",
    "1111111010000101",
    "1111101010111100",
    "1111010111100111",
    "1111000011001011",
    "1110110001100010",
    "1110100101101111",
    "1110100001000101",
    "1110100010111101",
    "1110101001001110",
    "1110110001011010",
    "1110111001101101",
    "1111000001010100",
    "1111001000011101",
    "1111001111101000",
    "1111010111101010",
    "1111100011100010",
    "1111110110101011",
    "1111101101110011",
    "1111001011111101",
    "1110101001000001",
    "1110001011101000",
    "1101111001011101",
    "1101110101111011",
    "1101111111111011",
    "1110010001100010",
    "1110100011100100",
    "1110101111111011",
    "1110110011110100",
    "1110110000100011",
    "1110101001011011",
    "1110100010011111",
    "1110100000101001",
    "1110101000101000",
    "1110111100111000",
    "1111011100010001",
    "1111111101111101",
    "1111011000111100",
    "1110111011010100",
    "1110101010000010",
    "1110100111010000",
    "1110110000110000",
    "1111000001000111",
    "1111010010001010",
    "1111011111001100",
    "1111100111101110",
    "1111101110111011",
    "1111111000101100",
    "1111111000010101",
    "1111100100111011",
    "1111010001001101",
    "1111000010011101",
    "1110111101001111",
    "1111000011100010",
    "1111010011010111",
    "1111101000001010",
    "1111111101001111",
    "1111110000101101",
    "1111100011001000",
    "1111011010011000",
    "1111010110100101",
    "1111010111110101",
    "1111011110100011",
    "1111101011011101",
    "1111111110100101",
    "1111101001011111",
    "1111010000000000",
    "1110111001010101",
    "1110101001011110",
    "1110100010100111",
    "1110100100010101",
    "1110101100100001",
    "1110111010000001",
    "1111001101101011",
    "1111101000101100",
    "1111110101001110",
    "1111001110110000",
    "1110101001010000",
    "1110001011000110",
    "1101111010000010",
    "1101111010001100",
    "1110001100100001",
    "1110101110110110",
    "1111011100011011",
    "1111110001011111",
    "1111000010001101",
    "1110011100000001",
    "1110000011011000",
    "1101111001100011",
    "1101111100001100",
    "1110000110111110",
    "1110010100101110",
    "1110100001010000",
    "1110101010010011",
    "1110110000011001",
    "1110111000001100",
    "1111000111111100",
    "1111100011010101",
    "1111110110101110",
    "1111001100100001",
    "1110100110101111",
    "1110001101010010",
    "1110000101100000",
    "1110010000010101",
    "1110101010011000",
    "1111001101111101",
    "1111110100101001",
    "1111100111100010",
    "1111001011000010",
    "1110111000101000",
    "1110110001010010",
    "1110110011111100",
    "1110111110100110",
    "1111001111110110",
    "1111100111100010",
    "1111111010010001",
    "1111010111010001",
    "1110110011010010",
    "1110010011010011",
    "1101111011101101",
    "1101101111011010",
    "1101101111001111",
    "1101111001011011",
    "1110001010001100",
    "1110011100110101",
    "1110101101010110",
    "1110111001101101",
    "1111000001111101",
    "1111000111101111",
    "1111001110101000",
    "1111011010101111",
    "1111101101111111",
    "1111111000110001",
    "1111011110000100",
    "1111001000011101",
    "1110111110001111",
    "1111000011111011",
    "1111011010111000",
    "1111111111110110",
    "1111010010101110",
    "1110100101110001",
    "1110000000110001",
    "1101101000111110",
    "1101100000010010",
    "1101100101110111",
    "1101110110001101",
    "1110001101010001",
    "1110101001010110",
    "1111001001110101",
    "1111101101101101",
    "1111101101011110",
    "1111001100001100",
    "1110110011011100",
    "1110100111000011",
    "1110101000001000",
    "1110110011100111",
    "1111000011011000",
    "1111010001001010",
    "1111011000101000",
    "1111011001110000",
    "1111011001000001",
    "1111011011111000",
    "1111100110010110",
    "1111111000111000",
    "1111110000011100",
    "1111011011100011",
    "1111001101101000",
    "1111001001010001",
    "1111001101001100",
    "1111010101010010",
    "1111011101001010",
    "1111100010010000",
    "1111100100100000",
    "1111100101101001",
    "1111100111101101",
    "1111101100100010",
    "1111110101000010",
    "1111111111010111",
    "1111110010010001",
    "1111100101101001",
    "1111011011010001",
    "1111010100010000",
    "1111010000101011",
    "1111001111111011",
    "1111010001010111",
    "1111010100101001",
    "1111011010010011",
    "1111100011100001",
    "1111110001001111",
    "1111111100011110",
    "1111100111100011",
    "1111010011001101",
    "1111000011001101",
    "1110111010110010",
    "1110111011011000",
    "1111000100101001",
    "1111010100111100",
    "1111101010000111",
    "1111111110010001",
    "1111100110101000",
    "1111010001000000",
    "1110111111001000",
    "1110110010011100",
    "1110101011111010",
    "1110101011111101",
    "1110110010110100",
    "1111000001010111",
    "1111011000010011",
    "1111110110101111",
    "1111100110101111",
    "1111000101101001",
    "1110101011110010",
    "1110011101111000",
    "1110011110011011",
    "1110101101001010",
    "1111000111000100",
    "1111100111010011",
    "1111110111011010",
    "1111011001100011",
    "1111000001110110",
    "1110110001101011",
    "1110101000111111",
    "1110100111010000",
    "1110101100111000",
    "1110111011011000",
    "1111010011100100",
    "1111110100010000",
    "1111100110010101",
    "1111000010000000",
    "1110100100011010",
    "1110010001110001",
    "1110001011011001",
    "1110001111011111",
    "1110011011001110",
    "1110101100100001",
    "1111000010011001",
    "1111011100010100",
    "1111111001000110",
    "1111101001010101",
    "1111001101110101",
    "1110110111101000",
    "1110101001101000",
    "1110100100101001",
    "1110100111101100",
    "1110110001011110",
    "1111000001001010",
    "1111010110110010",
    "1111110010001001",
    "1111101110000111",
    "1111001101001010",
    "1110101111011001",
    "1110011001011000",
    "1110001101111011",
    "1110001101000100",
    "1110010100100101",
    "1110100001010100",
    "1110110000100011",
    "1111000000111101",
    "1111010010100110",
    "1111100101111011",
    "1111111010110010",
    "1111101111111111",
    "1111011100011011",
    "1111001100100101",
    "1111000010010100",
    "1110111110101101",
    "1111000001111011",
    "1111001011101101",
    "1111011011101010",
    "1111110001100010",
    "1111110011001001",
    "1111010100010010",
    "1110110101000001",
    "1110011001101010",
    "1110000110100100",
    "1101111110110001",
    "1110000011000011",
    "1110010001010000",
    "1110100110001110",
    "1111000000010101",
    "1111011111010010",
    "1111111101010100",
    "1111010111001000",
    "1110110001110100",
    "1110010010011001",
    "1101111101101011",
    "1101110111000001",
    "1101111101110111",
    "1110001101101101",
    "1110100000011110",
    "1110110000011110",
    "1110111010011011",
    "1110111111101000",
    "1111000101101111",
    "1111010011000110",
    "1111101010110000",
    "1111110101100000",
    "1111010100011010",
    "1110111001101111",
    "1110101011101010",
    "1110101100010100",
    "1110111000000110",
    "1111001000001011",
    "1111010110001011",
    "1111011110010110",
    "1111100000001111",
    "1111011101101001",
    "1111011000110101",
    "1111010100001011",
    "1111010000111101",
    "1111001110110110",
    "1111001101010001",
    "1111001011010110",
    "1111001001100101",
    "1111001011000111",
    "1111010011101001",
    "1111100100101100",
    "1111111100011000",
    "1111101010001100",
    "1111010100101001",
    "1111000111000110",
    "1111000011100010",
    "1111001000100111",
    "1111010010011010",
    "1111011100011110",
    "1111100011000001",
    "1111100011110011",
    "1111011110001101",
    "1111010010100001",
    "1111000001111000",
    "1110101110101000",
    "1110011011100101",
    "1110001011111111",
    "1110000010100010",
    "1110000000101011",
    "1110000110011010",
    "1110010010001000",
    "1110100000110000",
    "1110101110110001",
    "1110111001101111",
    "1111000000111000",
    "1111000101111100",
    "1111001101000101",
    "1111011010010100",
    "1111101111011110",
    "1111110101000111",
    "1111011000011000",
    "1111000000000101",
    "1110110000111110",
    "1110101101100001",
    "1110110100100111",
    "1111000010010101",
    "1111010010010101",
    "1111100001001010",
    "1111101100111000",
    "1111110100100011",
    "1111110111101000",
    "1111110110000010",
    "1111110000011101",
    "1111100111111100",
    "1111011110010110",
    "1111010110011010",
    "1111010011011111",
    "1111011001001011",
    "1111101001010011",
    "1111111101000111",
    "1111011110001100",
    "1110111111100110",
    "1110100110100101",
    "1110010110110001",
    "1110010001001111",
    "1110010100101010",
    "1110011101111011",
    "1110101001110101",
    "1110110110100000",
    "1111000100011010",
    "1111010101001101",
    "1111101010001010",
    "1111111100111010",
    "1111100010011001",
    "1111001010000100",
    "1110110111101100",
    "1110101101100001",
    "1110101011010100",
    "1110101110011001",
    "1110110011010101",
    "1110110111110101",
    "1110111011110000",
    "1111000000010111",
    "1111000111000001",
    "1111010000010101",
    "1111011011111100",
    "1111101000010100",
    "1111110011011000",
    "1111111011010011",
    "1111111111010001",
    "1111111111111001",
    "1111111111000011",
    "1111111110111100",
    "1111111110110011",
    "1111111010000010",
    "1111110011111011",
    "1111101110100000",
    "1111101100000010",
    "1111101110010001",
    "1111110101110010",
    "1111111110000110",
    "1111101111001100",
    "1111011111111000",
    "1111010010101011",
    "1111001001101010",
    "1111000101111110",
    "1111000111100000",
    "1111001101100001",
    "1111010111101111",
    "1111100110010000",
    "1111111000111011",
    "1111110001011111",
    "1111011011110010",
    "1111001001001110",
    "1110111100101011",
    "1110110111111110",
    "1110111011010001",
    "1111000101010010",
    "1111010011101001",
    "1111100011110100",
    "1111110011100110",
    "1111111110101010",
    "1111110100110000",
    "1111110000001100",
    "1111110010001001",
    "1111111010110111",
    "1111110110101100",
    "1111100101001011",
    "1111010100001011",
    "1111000111100010",
    "1111000010000110",
    "1111000100101001",
    "1111001101100001",
    "1111011001001011",
    "1111100011100110",
    "1111101001110001",
    "1111101010001110",
    "1111100100110011",
    "1111011010010001",
    "1111001100000101",
    "1110111100011001",
    "1110101101110000",
    "1110100010111011",
    "1110011110011011",
    "1110100001111001",
    "1110101101011001",
    "1110111110111000",
    "1111010011010011",
    "1111101000100101",
    "1111111110010000",
    "1111101011001010",
    "1111010011101001",
    "1110111100010100",
    "1110100111100111",
    "1110011000110100",
    "1110010011000011",
    "1110010111011010",
    "1110100100000001",
    "1110110100110011",
    "1111000100111100",
    "1111010000111011",
    "1111011000010001",
    "1111011110011001",
    "1111101000011011",
    "1111111010001001",
    "1111101100010010",
    "1111001111001000",
    "1110110101000110",
    "1110100100111011",
    "1110100011010000",
    "1110110000010001",
    "1111000111111001",
    "1111100100000101",
    "1111111110101001",
    "1111101101000000",
    "1111100001100110",
    "1111011111111111",
    "1111100111010100",
    "1111110101001001",
    "1111111001011011",
    "1111100111111100",
    "1111011001110101",
    "1111010010000011",
    "1111010010101011",
    "1111011100010011",
    "1111101101011010",
    "1111111101011010",
    "1111101000100001",
    "1111010111011111",
    "1111001100010100",
    "1111000111010101",
    "1111000111011111",
    "1111001010110101",
    "1111001111011001",
    "1111010011010111",
    "1111010101010111",
    "1111010100100111",
    "1111010001001111",
    "1111001100001111",
    "1111000111011011",
    "1111000101000101",
    "1111000111011011",
    "1111010000000010",
    "1111011111001010",
    "1111110011111100",
    "1111110011110111",
    "1111011011100001",
    "1111000110010110",
    "1110110110111111",
    "1110101110101110",
    "1110101101100011",
    "1110110010011010",
    "1110111011100000",
    "1111000110111011",
    "1111010011011111",
    "1111100001001100",
    "1111110000100100",
    "1111111110010010",
    "1111101100010101",
    "1111011011100011",
    "1111001110100100",
    "1111000111101101",
    "1111001000011010",
    "1111010000111001",
    "1111100000010100",
    "1111110100110101",
    "1111110100001001",
    "1111011101110111",
    "1111001011011001",
    "1110111111001000",
    "1110111010001111",
    "1110111011110101",
    "1111000010010010",
    "1111001110000010",
    "1111100000011001",
    "1111111001011001",
    "1111101000110111",
    "1111001011001010",
    "1110110011001011",
    "1110100101100100",
    "1110100101000011",
    "1110110000010101",
    "1111000010011111",
    "1111010101100010",
    "1111100101110001",
    "1111110100100010",
    "1111111010000110",
    "1111100011110110",
    "1111001001001100",
    "1110101110010100",
    "1110011001101011",
    "1110010001000101",
    "1110010111010110",
    "1110101010000111",
    "1111000010100110",
    "1111011001011110",
    "1111101001100000",
    "1111110001101101",
    "1111110100101001",
    "1111110101010111",
    "1111111000001010",
    "1111111101111001",
    "1111101010011111",
    "1111001110100011",
    "1110101110101000",
    "1110010001101110",
    "1101111110001101",
    "1101111000001100",
    "1110000000011010",
    "1110010011011010",
    "1110101011001110",
    "1111000001101011",
    "1111010001101100",
    "1111011010000110",
    "1111011110101001",
    "1111100101011010",
    "1111110011100001",
    "1111110101011010",
    "1111011000111110",
    "1110111101100100",
    "1110101010001001",
    "1110100011110100",
    "1110101010110111",
    "1110111010011011",
    "1111001011101101",
    "1111011001000001",
    "1111011111101011",
    "1111100000101110",
    "1111100000011010",
    "1111100100110100",
    "1111110010100100",
    "1111110101110111",
    "1111011000110000",
    "1110111100111000",
    "1110101000101100",
    "1110011111011100",
    "1110100000000010",
    "1110100101110111",
    "1110101011011101",
    "1110101100101101",
    "1110100111111111",
    "1110011110101101",
    "1110010100000011",
    "1110001011111101",
    "1110001001010001",
    "1110001100111000",
    "1110010101101010",
    "1110100001000111",
    "1110101100010111",
    "1110110101100000",
    "1110111101011100",
    "1111001000100000",
    "1111011011000001",
    "1111110110010110",
    "1111100111111100",
    "1111000101110001",
    "1110101001010011",
    "1110010111011011",
    "1110010010001010",
    "1110010110111001",
    "1110011111111111",
    "1110101000000011",
    "1110101100111100",
    "1110110001010010",
    "1110111001101101",
    "1111001001011110",
    "1111100001000111",
    "1111111101100011",
    "1111100110100001",
    "1111010000011110",
    "1111000011001011",
    "1110111110010010",
    "1110111110111101",
    "1111000001101110",
    "1111000100011000",
    "1111000111000011",
    "1111001011011001",
    "1111010011010000",
    "1111011111010001",
    "1111101110011110",
    "1111111110010000",
    "1111110100110110",
    "1111101110001110",
    "1111101111101000",
    "1111111000101100",
    "1111111000101111",
    "1111100111101110",
    "1111010111011000",
    "1111001010011110",
    "1111000011000110",
    "1111000010000000",
    "1111000110110100",
    "1111010000011100",
    "1111011101111010",
    "1111101110101110",
    "1111111100111001",
    "1111100100100100",
    "1111001000010011",
    "1110101001101000",
    "1110001011111000",
    "1101110011101110",
    "1101100101101010",
    "1101100100010111",
    "1101101111011100",
    "1110000011101110",
    "1110011011111000",
    "1110110011111011",
    "1111001100010100",
    "1111100111111011",
    "1111110110111100",
    "1111010000011111",
    "1110101000110111",
    "1110000110100000",
    "1101110000001100",
    "1101101010101000",
    "1101110101000110",
    "1110001010001110",
    "1110100011000011",
    "1110111010111010",
    "1111010010100010",
    "1111101101010000",
    "1111110010111100",
    "1111001110100110",
    "1110101001110010",
    "1110001011000111",
    "1101111000101000",
    "1101110101100100",
    "1101111111111101",
    "1110010001110110",
    "1110100101010010",
    "1110110110110111",
    "1111000110110110",
    "1111010111001001",
    "1111101000011011",
    "1111111001100101",
    "1111110111111101",
    "1111101111001010",
    "1111101101010011",
    "1111110001001011",
    "1111110111100101",
    "1111111100101110",
    "1111111101110001",
    "1111111010011001",
    "1111110100100101",
    "1111101111000101",
    "1111101011110111",
    "1111101011001100",
    "1111101100000111",
    "1111101101010010",
    "1111101101010010",
    "1111101011010000",
    "1111100110111011",
    "1111100000011010",
    "1111010111101100",
    "1111001100100011",
    "1110111111000100",
    "1110110000100111",
    "1110100011111001",
    "1110011011111000",
    "1110011011000010",
    "1110100010001000",
    "1110110000010111",
    "1111000100001011",
    "1111011011101111",
    "1111110101011101",
    "1111101111110100",
    "1111010101000001",
    "1110111011000010",
    "1110100011101001",
    "1110010001011100",
    "1110000110110001",
    "1110000100100000",
    "1110001001101000",
    "1110010011011101",
    "1110011111000101",
    "1110101001101011",
    "1110110010101111",
    "1110111101011100",
    "1111001110010010",
    "1111100111111101",
    "1111110110101001",
    "1111010010101111",
    "1110110011001111",
    "1110011110001111",
    "1110010111010101",
    "1110011101011110",
    "1110101100000111",
    "1110111101100011",
    "1111001100110101",
    "1111010111011111",
    "1111011101100000",
    "1111011111111101",
    "1111100000011111",
    "1111100000011111",
    "1111100000000011",
    "1111011111001000",
    "1111011101101000",
    "1111011011011110",
    "1111011001001011",
    "1111010111011101",
    "1111010110110111",
    "1111010111011011",
    "1111011000101010",
    "1111011010010100",
    "1111011100100000",
    "1111100000000010",
    "1111100111100001",
    "1111110101111111",
    "1111110011001100",
    "1111010101011101",
    "1110110101000001",
    "1110010111101101",
    "1110000011000001",
    "1101111010101000",
    "1101111110100011",
    "1110001011011011",
    "1110011100010110",
    "1110101100101000",
    "1110111001010000",
    "1111000001100110",
    "1111000110011000",
    "1111001001000001",
    "1111001100110111",
    "1111010110010000",
    "1111100111101100",
    "1111111111100010",
    "1111100011111100",
    "1111001100001100",
    "1110111110001010",
    "1110111101100011",
    "1111001010100011",
    "1111100000100111",
    "1111111000111111",
    "1111110010011011",
    "1111100101000110",
    "1111011110110000",
    "1111011101011100",
    "1111011111101001",
    "1111100100100100",
    "1111101100100111",
    "1111111000100101",
    "1111110111110101",
    "1111100110011101",
    "1111010110000100",
    "1111001001111101",
    "1111000100001011",
    "1111000100101111",
    "1111001001101010",
    "1111010000001010",
    "1111011000010001",
    "1111100100110111",
    "1111111000010101",
    "1111101101000101",
    "1111001110001111",
    "1110110000100100",
    "1110011001110010",
    "1110001110011100",
    "1110010000000000",
    "1110011011000111",
    "1110101001110100",
    "1110110111000100",
    "1111000001111011",
    "1111001101101000",
    "1111011101101011",
    "1111110010111111",
    "1111110100111110",
    "1111100000010010",
    "1111010110010000",
    "1111011100011100",
    "1111110011110100",
    "1111101000001110",
    "1110111111111010",
    "1110011011011101",
    "1110000000011001",
    "1101110000010100",
    "1101101010000100",
    "1101101011001111",
    "1101110001001010",
    "1101111001110000",
    "1110000011111000",
    "1110001110110000",
    "1110011001111010",
    "1110100100100010",
    "1110101101101001",
    "1110110100111001",
    "1110111011001100",
    "1111000010011001",
    "1111001100101000",
    "1111011011011000",
    "1111101110111001",
    "1111111001111111",
    "1111100010000010",
    "1111001100110000",
    "1110111101000101",
    "1110110100011010",
    "1110110010011001",
    "1110110101010000",
    "1110111010110000",
    "1111000000101011",
    "1111000100111110",
    "1111000110011101",
    "1111000100101100",
    "1111000000010111",
    "1110111011101111",
    "1110111001101011",
    "1110111100110000",
    "1111000110001011",
    "1111010100111011",
    "1111100101110110",
    "1111110100011000",
    "1111111100010000",
    "1111111011001111",
    "1111110001111001",
    "1111100011001000",
    "1111010011001111",
    "1111000110011000",
    "1110111111111010",
    "1111000001111110",
    "1111001101001111",
    "1111100000101110",
    "1111111010011001",
    "1111101000101101",
    "1111001100010110",
    "1110110100001101",
    "1110100011011100",
    "1110011011111100",
    "1110011101111111",
    "1110101000110111",
    "1110111011100011",
    "1111010100100101",
    "1111110001110110",
    "1111101111101111",
    "1111010011111100",
    "1110111110001101",
    "1110110000110101",
    "1110101100000010",
    "1110101101111000",
    "1110110011001011",
    "1110111000111010",
    "1110111101011110",
    "1111000001000011",
    "1111000101001001",
    "1111001011110010",
    "1111010110010110",
    "1111100100111110",
    "1111110110010111",
    "1111110111101001",
    "1111100111100010",
    "1111011011010100",
    "1111010100010101",
    "1111010011001011",
    "1111010111110111",
    "1111100001111110",
    "1111110000110000",
    "1111111101000110",
    "1111101001101010",
    "1111010111011101",
    "1111001001010101",
    "1111000001110100",
    "1111000010100100",
    "1111001011101000",
    "1111011011100000",
    "1111101111010010",
    "1111111100011011",
    "1111101010101001",
    "1111011100110111",
    "1111010011010101",
    "1111001101100011",
    "1111001010111010",
    "1111001011001010",
    "1111001110010111",
    "1111010101011101",
    "1111100010100010",
    "1111110111011000",
    "1111101100000111",
    "1111001010101000",
    "1110101000111100",
    "1110001100110010",
    "1101111011000010",
    "1101110110001101",
    "1101111101011001",
    "1110001100110000",
    "1110011111101001",
    "1110110100011111",
    "1111001100110000",
    "1111101010001010",
    "1111110011101001",
    "1111010000010001",
    "1110110001011001",
    "1110011100111101",
    "1110010111001101",
    "1110100000001010",
    "1110110011001101",
    "1111001001100000",
    "1111011100101011",
    "1111101000111011",
    "1111101110001011",
    "1111101110010010",
    "1111101011100011",
    "1111100111111101",
    "1111100100000011",
    "1111011111111010",
    "1111011101110000",
    "1111100001110001",
    "1111101111100011",
    "1111110111110001",
    "1111010111010011",
    "1110110101101001",
    "1110011010100010",
    "1110001011111101",
    "1110001011011011",
    "1110010100111011",
    "1110100010000011",
    "1110101100110010",
    "1110110001011001",
    "1110110001100001",
    "1110110011001101",
    "1110111100101010",
    "1111010001000010",
    "1111101110010010",
    "1111110010010011",
    "1111011000010011",
    "1111001001011110",
    "1111001000001001",
    "1111010010010000",
    "1111100100010111",
    "1111111011011100",
    "1111101010101101",
    "1111001111101011",
    "1110110101100100",
    "1110011111101001",
    "1110010000111110",
    "1110001011101011",
    "1110001111111111",
    "1110011100010001",
    "1110101111010110",
    "1111001000011010",
    "1111100110001000",
    "1111111001111001",
    "1111011011011011",
    "1111000010011101",
    "1110110010100110",
    "1110101110100100",
    "1110110110100100",
    "1111000111011010",
    "1111011100000101",
    "1111110001000001",
    "1111111010010011",
    "1111100100100100",
    "1111001100100000",
    "1110110010101100",
    "1110011010001011",
    "1110000111011111",
    "1101111111010010",
    "1110000100001011",
    "1110010101010010",
    "1110101110100001",
    "1111001010101111",
    "1111100101010011",
    "1111111011011011",
    "1111110100010101",
    "1111101010011001",
    "1111100101111100",
    "1111100101101111",
    "1111101000100010",
    "1111101101010000",
    "1111110011000101",
    "1111111001010000",
    "1111111110110100",
    "1111111101000100",
    "1111111010110101",
    "1111111010001000",
    "1111111010100110",
    "1111111100010001",
    "1111111111011111",
    "1111111011101110",
    "1111110101111011",
    "1111101111111100",
    "1111101010101000",
    "1111100111000110",
    "1111100110100110",
    "1111101010000100",
    "1111110001111000",
    "1111111101110100",
    "1111110010101100",
    "1111100001000010",
    "1111001110111111",
    "1110111110110000",
    "1110110010001010",
    "1110101010011001",
    "1110100111111010",
    "1110101010100000",
    "1110110001001000",
    "1110111010001100",
    "1111000011111110",
    "1111001100111100",
    "1111010100011100",
    "1111011010101101",
    "1111100000000000",
    "1111100101100101",
    "1111101110110011",
    "1111111110101001",
    "1111101010010110",
    "1111001110111000",
    "1110110100100000",
    "1110100001010111",
    "1110011001100010",
    "1110011110110011",
    "1110110000110001",
    "1111001100111111",
    "1111101111010111",
    "1111101101011000",
    "1111001110110000",
    "1110111000111111",
    "1110101111000010",
    "1110110001110110",
    "1110111111010110",
    "1111010011001010",
    "1111101001101101",
    "1111111101111001",
    "1111100011000110",
    "1111000101100101",
    "1110100111011010",
    "1110001100010111",
    "1101111000001011",
    "1101101101111111",
    "1101101111011110",
    "1101111010101011",
    "1110001011001110",
    "1110011011101010",
    "1110100111100000",
    "1110101100111010",
    "1110101100111000",
    "1110101010001001",
    "1110100111100101",
    "1110100111100101",
    "1110101101000100",
    "1110111010111100",
    "1111010001011100",
    "1111101101111000",
    "1111110101000000",
    "1111011101101110",
    "1111010001100001",
    "1111010011010101",
    "1111100001110000",
    "1111110110100101",
    "1111110100001110",
    "1111100000110011",
    "1111001101110101",
    "1110111001010001",
    "1110100010111101",
    "1110001101110010",
    "1101111110000010",
    "1101111000000100",
    "1101111110100110",
    "1110010000000000",
    "1110100110111001",
    "1110111100101110",
    "1111001011101011",
    "1111010010010000",
    "1111010101101010",
    "1111011101101000",
    "1111101111110111",
    "1111110010111011",
    "1111010000100100",
    "1110110001110110",
    "1110011110111010",
    "1110011101010100",
    "1110101100110101",
    "1111001000001110",
    "1111101000111000",
    "1111110111000111",
    "1111011011111000",
    "1111000111101111",
    "1110111101000100",
    "1110111101101101",
    "1111001001111100",
    "1111100000111001",
    "1111111111110101",
    "1111011101111101",
    "1110111110001101",
    "1110100110100000",
    "1110011010011001",
    "1110011001111001",
    "1110100001101110",
    "1110101101010110",
    "1110111001001001",
    "1111000101000110",
    "1111010100100100",
    "1111101010101000",
    "1111110111111101",
    "1111010110010000",
    "1110110101111110",
    "1110011100100001",
    "1110001101110000",
    "1110001010010011",
    "1110001111001100",
    "1110011001010000",
    "1110100111100111",
    "1110111010110100",
    "1111010011111001",
    "1111110010011010",
    "1111101100011110",
    "1111001100110011",
    "1110110011010011",
    "1110100011111001",
    "1110011111001100",
    "1110100011011010",
    "1110101110001101",
    "1110111110000111",
    "1111010010111011",
    "1111101100111011",
    "1111110100100010",
    "1111010100000001",
    "1110110110000011",
    "1110011111111011",
    "1110010101100000",
    "1110010111110100",
    "1110100100101010",
    "1110110111010110",
    "1111001010010110",
    "1111011001010011",
    "1111100011110011",
    "1111101101010110",
    "1111111010010100",
    "1111110010111110",
    "1111011011110111",
    "1111000100111001",
    "1110110011101001",
    "1110101100110101",
    "1110110010010010",
    "1111000001011010",
    "1111010101010011",
    "1111101010011100",
    "1111111111111100",
    "1111101001101101",
    "1111010010100100",
    "1110111100100110",
    "1110101011010001",
    "1110100010101001",
    "1110100111001001",
    "1110111011101000",
    "1111011111001010",
    "1111110011001011",
    "1111000011010010",
    "1110011001101000",
    "1101111100110111",
    "1101110000010010",
    "1101110011100010",
    "1110000010110011",
    "1110011000100010",
    "1110101111010100",
    "1111000010111000",
    "1111010010101100",
    "1111100010101110",
    "1111110111100110",
    "1111101100001010",
    "1111001001111001",
    "1110100110101101",
    "1110001001010001",
    "1101110111111100",
    "1101110110001011",
    "1110000001110011",
    "1110010100110111",
    "1110101000110010",
    "1110111000110100",
    "1111000011011100",
    "1111001001011011",
    "1111001100010110",
    "1111001110100001",
    "1111010001100001",
    "1111010110110111",
    "1111100001010010",
    "1111110010100010",
    "1111110101110010",
    "1111011010010011",
    "1110111111101001",
    "1110101010110111",
    "1110100000000010",
    "1110100000111000",
    "1110101010110101",
    "1110111000101100",
    "1111000110010110",
    "1111010010001111",
    "1111011100110011",
    "1111100110111110",
    "1111101111111111",
    "1111110101101011",
    "1111110101000000",
    "1111101011000000",
    "1111010111011111",
    "1110111110001010",
    "1110100101010011",
    "1110010011011100",
    "1110001100101011",
    "1110010001001100",
    "1110011101110011",
    "1110101101101101",
    "1110111100100110",
    "1111001001010101",
    "1111010110011010",
    "1111100111110001",
    "1111111111110110",
    "1111100010100111",
    "1111000100100101",
    "1110101100010110",
    "1110011111001111",
    "1110011111011110",
    "1110101011011011",
    "1110111111011001",
    "1111010111011000",
    "1111110000010010",
    "1111110111100101",
    "1111100001001010",
    "1111001101100000",
    "1110111110001101",
    "1110110101110110",
    "1110110110111110",
    "1111000010111001",
    "1111011000111111",
    "1111110110111001",
    "1111100111011010",
    "1111000110110111",
    "1110101011111000",
    "1110011001010110",
    "1110001111111010",
    "1110001110100001",
    "1110010010111000",
    "1110011010011000",
    "1110100100101001",
    "1110110011100110",
    "1111001000101101",
    "1111100011110001",
    "1111111101110111",
    "1111100000111101",
    "1111001010010110",
    "1110111110000101",
    "1110111101010100",
    "1111000101010000",
    "1111010001001111",
    "1111011101011110",
    "1111101001000100",
    "1111110101111101",
    "1111111001100111",
    "1111100100111001",
    "1111001101011001",
    "1110110111000011",
    "1110100111000011",
    "1110100001011111",
    "1110100111111111",
    "1110111000110101",
    "1111010000001100",
    "1111101010000101",
    "1111111011111010",
    "1111100010010000",
    "1111001000100011",
    "1110101111000111",
    "1110010111101100",
    "1110000101001101",
    "1101111010101000",
    "1101111001110010",
    "1110000010100111",
    "1110010011000110",
    "1110100111111001",
    "1110111101101101",
    "1111010011110011",
    "1111101100000010",
    "1111110111100001",
    "1111010110110111",
    "1110110100110111",
    "1110010110101111",
    "1110000010000101",
    "1101111010111010",
    "1110000001101001",
    "1110010010010111",
    "1110100110111100",
    "1110111001100000",
    "1111000110111111",
    "1111010001011010",
    "1111011101110000",
    "1111110000010001",
    "1111110110001000",
    "1111011001000111",
    "1110111111010100",
    "1110101111100001",
    "1110101110011110",
    "1110111100100000",
    "1111010100110100",
    "1111110000001011",
    "1111111000000111",
    "1111101000010110",
    "1111100001111110",
    "1111100100110110",
    "1111101111100100",
    "1111111111110001",
    "1111101101000101",
    "1111011001100101",
    "1111001000001100",
    "1110111011011011",
    "1110110101011000",
    "1110110111011000",
    "1111000001000111",
    "1111010000011001",
    "1111100001101110",
    "1111110001011101",
    "1111111100111010",
    "1111111101010001",
    "1111111101000100",
    "1111111111000101",
    "1111111001100011",
    "1111110100110101",
    "1111110011001001",
    "1111110110001110",
    "1111111110111101",
    "1111110010110110",
    "1111100000101011",
    "1111001101000100",
    "1110111011010110",
    "1110101110101000",
    "1110101001000111",
    "1110101011101011",
    "1110110101101110",
    "1111000101100100",
    "1111011001101111",
    "1111110001011110",
    "1111110011110011",
    "1111010111011011",
    "1110111100000100",
    "1110100101001011",
    "1110010101101100",
    "1110001111010001",
    "1110010001010010",
    "1110011001010001",
    "1110100011111011",
    "1110101110110011",
    "1110111001011101",
    "1111000101001110",
    "1111010011110011",
    "1111100110000100",
    "1111111011100000",
    "1111101110000010",
    "1111011001011011",
    "1111001001000110",
    "1110111110011110",
    "1110111001101101",
    "1110111001110101",
    "1110111101011110",
    "1111000011000011",
    "1111001001001100",
    "1111001110110011",
    "1111010010110110",
    "1111010101000001",
    "1111010101110110",
    "1111010110010110",
    "1111010111101111",
    "1111011010101010",
    "1111011111000000",
    "1111100100011000",
    "1111101010011100",
    "1111110001011011",
    "1111111010001111",
    "1111111010000111",
    "1111101011010011",
    "1111011001110000",
    "1111000111001110",
    "1110110110001001",
    "1110101000111111",
    "1110100001010100",
    "1110011111011001",
    "1110100001111000",
    "1110100110100000",
    "1110101010101000",
    "1110101100010100",
    "1110101011000100",
    "1110100111111010",
    "1110100100111110",
    "1110100100100010",
    "1110101000001011",
    "1110110000000111",
    "1110111011100101",
    "1111001001100011",
    "1111011001111001",
    "1111101101000101",
    "1111111100101001",
    "1111100100010011",
    "1111001100011110",
    "1110111000101100",
    "1110101100011100",
    "1110101001110101",
    "1110110000010100",
    "1110111101000010",
    "1111001011110010",
    "1111011000100101",
    "1111100000110000",
    "1111100011011100",
    "1111100001011001",
    "1111011101001110",
    "1111011011100011",
    "1111100000110101",
    "1111101111000101",
    "1111111010111010",
    "1111100001100111",
    "1111001010110000",
    "1110111011001100",
    "1110110101100000",
    "1110111000100111",
    "1111000000001100",
    "1111000110111001",
    "1111001000100011",
    "1111000100000101",
    "1110111011101000",
    "1110110010111110",
    "1110101101110000",
    "1110101110000111",
    "1110110011101111",
    "1110111100100001",
    "1111000101101100",
    "1111001101000000",
    "1111010001110001",
    "1111010101001000",
    "1111011011001100",
    "1111101001001001",
    "1111111110011001",
    "1111011100101010",
    "1110110110101111",
    "1110010100010101",
    "1101111100011011",
    "1101110011100111",
    "1101111001111100",
    "1110001010011000",
    "1110011110001001",
    "1110101111011100",
    "1110111011001010",
    "1111000010011001",
    "1111001001011011",
    "1111010101100000",
    "1111101010011000",
    "1111111000011000",
    "1111010111010101",
    "1110111000101111",
    "1110100010101001",
    "1110011000110100",
    "1110011010111100",
    "1110100101100101",
    "1110110100010010",
    "1111000011010101",
    "1111010000110001",
    "1111011100000010",
    "1111100101001101",
    "1111101100101110",
    "1111110010101011",
    "1111110111101000",
    "1111111101111110",
    "1111110111110011",
    "1111101000110101",
    "1111010110001011",
    "1111000011000101",
    "1110110011100110",
    "1110101011011101",
    "1110101100110111",
    "1110110110101111",
    "1111000101001110",
    "1111010011111110",
    "1111011111100110",
    "1111100111001100",
    "1111101011110001",
    "1111101110101111",
    "1111110001010000",
    "1111110011110011",
    "1111110101110101",
    "1111110110110001",
    "1111110110011000",
    "1111110100111010",
    "1111110011010010",
    "1111110010100010",
    "1111110011010000",
    "1111110101100001",
    "1111111001001110",
    "1111111110101000",
    "1111111001011010",
    "1111101110010100",
    "1111100000011100",
    "1111010001010100",
    "1111000011101110",
    "1110111010100011",
    "1110110111110111",
    "1110111100001100",
    "1111000110010011",
    "1111010011100001",
    "1111100000111000",
    "1111101100010011",
    "1111110101001000",
    "1111111100000111",
    "1111111100011101",
    "1111110001000100",
    "1111011110110110",
    "1111000101101100",
    "1110101000011010",
    "1110001011110000",
    "1101110100110111",
    "1101100111100111",
    "1101100101101110",
    "1101101110000100",
    "1101111101010100",
    "1110001111100100",
    "1110100001010000",
    "1110110000111101",
    "1111000000001101",
    "1111010010010000",
    "1111101001100010",
    "1111111010000110",
    "1111011100010001",
    "1111000010101001",
    "1110110010111011",
    "1110110001001000",
    "1110111101011011",
    "1111010100010011",
    "1111110000011110",
    "1111110011010001",
    "1111011010011110",
    "1111000110100000",
    "1110110111100111",
    "1110101101000010",
    "1110100110000000",
    "1110100010011111",
    "1110100010111101",
    "1110100111110111",
    "1110110001011001",
    "1110111110110000",
    "1111001110000111",
    "1111011101000010",
    "1111101000110111",
    "1111101110111111",
    "1111101101001101",
    "1111100010010000",
    "1111001111001100",
    "1110110111100010",
    "1110100000100001",
    "1110001111100001",
    "1110001000001001",
    "1110001011000001",
    "1110010101111001",
    "1110100100110110",
    "1110110101100010",
    "1111001001011011",
    "1111100011000110",
    "1111111100000110",
    "1111010101110110",
    "1110101111001101",
    "1110001110101000",
    "1101111001111010",
    "1101110100011000",
    "1101111100001110",
    "1110001011110010",
    "1110011100101110",
    "1110101011001110",
    "1110111001000001",
    "1111001010110100",
    "1111100011111110",
    "1111111010111111",
    "1111010110001101",
    "1110110100101111",
    "1110011101011100",
    "1110010100011100",
    "1110011000111110",
    "1110100101111001",
    "1110110100110011",
    "1111000000101001",
    "1111000111100010",
    "1111001010100110",
    "1111001011101011",
    "1111001100101110",
    "1111010001001000",
    "1111011100100011",
    "1111110000101101",
    "1111110011100000",
    "1111010100011101",
    "1110111000000011",
    "1110100011010000",
    "1110011001100101",
    "1110011011101010",
    "1110100101101110",
    "1110110001111001",
    "1110111010100010",
    "1110111101001100",
    "1110111100111010",
    "1110111110110101",
    "1111000110111110",
    "1111010110011111",
    "1111101010000000",
    "1111111011011111",
    "1111111011000011",
    "1111111101110101",
    "1111110011101001",
    "1111011110010010",
    "1111001000011011",
    "1110110111100000",
    "1110101101110111",
    "1110101011000110",
    "1110101101100110",
    "1110110011001111",
    "1110111010000100",
    "1111000001101011",
    "1111001011011011",
    "1111011001110010",
    "1111101110010110",
    "1111110111101010",
    "1111011011101101",
    "1111000010001101",
    "1110101111001010",
    "1110100101001110",
    "1110100101011011",
    "1110101110100001",
    "1110111101010111",
    "1111001110000101",
    "1111011101101101",
    "1111101010101100",
    "1111110100111101",
    "1111111101010000",
    "1111111011001011",
    "1111110010101100",
    "1111100111101001",
    "1111011010000110",
    "1111001100000010",
    "1111000000111001",
    "1110111100000100",
    "1110111111011100",
    "1111001011001001",
    "1111011101000100",
    "1111110000111110",
    "1111111101110011",
    "1111110010101101",
    "1111101110100111",
    "1111110000000111",
    "1111110101001010",
    "1111111100001101",
    "1111111011010100",
    "1111110001010011",
    "1111100101001101",
    "1111010111001011",
    "1111001000100010",
    "1110111011111100",
    "1110110101000001",
    "1110110111011011",
    "1111000100111011",
    "1111011100011100",
    "1111111010001111",
    "1111100110111011",
    "1111001100011011",
    "1110111010001001",
    "1110110001111101",
    "1110110011000000",
    "1110111010101111",
    "1111000110000100",
    "1111010010010101",
    "1111011111010001",
    "1111101111101011",
    "1111111001010000",
    "1111011010101111",
    "1110110111001101",
    "1110010100010101",
    "1101111000101010",
    "1101101001100000",
    "1101101001001011",
    "1101110101011000",
    "1110001000101111",
    "1110011101101101",
    "1110110000000011",
    "1110111111010111",
    "1111001111100110",
    "1111100101001101",
    "1111111101101101",
    "1111011011010110",
    "1110111010001110",
    "1110100001111001",
    "1110010111111110",
    "1110011111000101",
    "1110110110100100",
    "1111011010110101",
    "1111111001100110",
    "1111001101010110",
    "1110100110100111",
    "1110001010101010",
    "1101111101001001",
    "1101111110111011",
    "1110001101001100",
    "1110100010000011",
    "1110110111100111",
    "1111001011100101",
    "1111011111110110",
    "1111110111010011",
    "1111101101000001",
    "1111001110111111",
    "1110110010100110",
    "1110011101001010",
    "1110010011110110",
    "1110011000010110",
    "1110100111110010",
    "1110111100010111",
    "1111010000010101",
    "1111100000110110",
    "1111101111011011",
    "1111111111110001",
    "1111101011000101",
    "1111010000111000",
    "1110110101001000",
    "1110011101011011",
    "1110001110111010",
    "1110001100010111",
    "1110010100111100",
    "1110100100111100",
    "1110110111110001",
    "1111001001101101",
    "1111011000111111",
    "1111100100111011",
    "1111101101110011",
    "1111110110010100",
    "1111111101011001",
    "1111101010111110",
    "1111010010111001",
    "1110111000111100",
    "1110100010100100",
    "1110010100100010",
    "1110010001110110",
    "1110011010100110",
    "1110101011000100",
    "1110111101100000",
    "1111001100010111",
    "1111010100001110",
    "1111010101101010",
    "1111010101100111",
    "1111011010110101",
    "1111101010010010",
    "1111111011110001",
    "1111011100100110",
    "1111000000000111",
    "1110101110000010",
    "1110101011001100",
    "1110110110100000",
    "1111001001101111",
    "1111011101001010",
    "1111101010101100",
    "1111101111101110",
    "1111101101000110",
    "1111100101010111",
    "1111011100000001",
    "1111010100001011",
    "1111001110111000",
    "1111001011011101",
    "1111001000101000",
    "1111000101100100",
    "1111000010010111",
    "1110111111101110",
    "1110111110010110",
    "1110111110010111",
    "1111000000110110",
    "1111001000100101",
    "1111011000011101",
    "1111110001011001",
    "1111101110011010",
    "1111001011100110",
    "1110101011110111",
    "1110010100000110",
    "1110000111001011",
    "1110000100010111",
    "1110001000111111",
    "1110010011010010",
    "1110100010111110",
    "1110111000011110",
    "1111010011010011",
    "1111110000110010",
    "1111110010111001",
    "1111011011110101",
    "1111001101010100",
    "1111001000100010",
    "1111001011111111",
    "1111010101001001",
    "1111100010000000",
    "1111110010001010",
    "1111111001100000",
    "1111100000100111",
    "1111000100001011",
    "1110100111011101",
    "1110001111010110",
    "1110000000011100",
    "1101111101010001",
    "1110000101001110",
    "1110010100111100",
    "1110100111110101",
    "1110111001110000",
    "1111001000011000",
    "1111010100011000",
    "1111100001000111",
    "1111110001100010",
    "1111111001110101",
    "1111100011111000",
    "1111010001110000",
    "1111001000110100",
    "1111001100111111",
    "1111011111000111",
    "1111111100011010",
    "1111100000001000",
    "1110111011110010",
    "1110011010110000",
    "1110000000001101",
    "1101101110010001",
    "1101100110010101",
    "1101101000101000",
    "1101110100001010",
    "1110000111110001",
    "1110100011010010",
    "1111000110011111",
    "1111101111100101",
    "1111100101010011",
    "1110111101110011",
    "1110011111001101",
    "1110001101100001",
    "1110001010100101",
    "1110010100110110",
    "1110100111110100",
    "1110111110000010",
    "1111010011111011",
    "1111101000111011",
    "1111111110001111",
    "1111101011010011",
    "1111010100100100",
    "1111000000010001",
    "1110110010100010",
    "1110101111101000",
    "1110111001011011",
    "1111001110011111",
    "1111101010000111",
    "1111111001111110",
    "1111100011101010",
    "1111010110101100",
    "1111010100010101",
    "1111011100000010",
    "1111101011100110",
    "1111111111110100",
    "1111101010110100",
    "1111010111101010",
    "1111001001001011",
    "1111000000111000",
    "1110111111101110",
    "1111000110001101",
    "1111010011101110",
    "1111100110010101",
    "1111111010101110",
    "1111110010101101",
    "1111100101011010",
    "1111011111101001",
    "1111100010001111",
    "1111101100001101",
    "1111111011000000",
    "1111110100101101",
    "1111100110011011",
    "1111011100110101",
    "1111011010000001",
    "1111011111001010",
    "1111101100010011",
    "1111111111101010",
    "1111101001110100",
    "1111010100000101",
    "1111000010100001",
    "1110110111010000",
    "1110110010101111",
    "1110110011101010",
    "1110110111110111",
    "1110111101010110",
    "1111000011010010",
    "1111001010010100",
    "1111010011011111",
    "1111011111001111",
    "1111101101000001",
    "1111111011011001",
    "1111110111100000",
    "1111101101011100",
    "1111100111101010",
    "1111100110111000",
    "1111101011001100",
    "1111110100010101",
    "1111111110000101",
    "1111101100100001",
    "1111010111111010",
    "1111000010000110",
    "1110101101110011",
    "1110011101111000",
    "1110010100100100",
    "1110010010111000",
    "1110011000100000",
    "1110100011101110",
    "1110110010110110",
    "1111000101110110",
    "1111011101010001",
    "1111111001000101",
    "1111101000011100",
    "1111001010111010",
    "1110110010011100",
    "1110100010100100",
    "1110011101010010",
    "1110100001110110",
    "1110101101010001",
    "1110111011111111",
    "1111001011010011",
    "1111011001111101",
    "1111100111111010",
    "1111110101001001",
    "1111111110100111",
    "1111110100100011",
    "1111101110100000",
    "1111101110010000",
    "1111110100110001",
    "1111111110000000",
    "1111101011011101",
    "1111010101101111",
    "1110111111010010",
    "1110101010101101",
    "1110011010100101",
    "1110010001100001",
    "1110010001110001",
    "1110011100110010",
    "1110110010100111",
    "1111010001111000",
    "1111110111100001",
    "1111100000110001",
    "1110111011111000",
    "1110011110010001",
    "1110001010111100",
    "1110000010110011",
    "1110000100100010",
    "1110001101010111",
    "1110011010000010",
    "1110100111110100",
    "1110110101000000",
    "1111000001000000",
    "1111001011111000",
    "1111010101110010",
    "1111011110101011",
    "1111100110100001",
    "1111101101011011",
    "1111110011010101",
    "1111110111101101",
    "1111111001100011",
    "1111110111101100",
    "1111110001010100",
    "1111100110100010",
    "1111011000101010",
    "1111001010000111",
    "1110111101111101",
    "1110110110111001",
    "1110110110100100",
    "1110111101000111",
    "1111001001111100",
    "1111011100011001",
    "1111110011111001",
    "1111110000101101",
    "1111010011110001",
    "1110111000100101",
    "1110100010101001",
    "1110010100101111",
    "1110010000001000",
    "1110010100000011",
    "1110011101111000",
    "1110101010000111",
    "1110110101100100",
    "1110111110001010",
    "1111000011001011",
    "1111000100111110",
    "1111000100100010",
    "1111000011001010",
    "1111000001110100",
    "1111000000111110",
    "1111000000100111",
    "1111000000010001",
    "1110111111111101",
    "1111000010010100",
    "1111001011010100",
    "1111011101000101",
    "1111110110110011",
    "1111101011110010",
    "1111010001000000",
    "1110111110100001",
    "1110111000000100",
    "1110111101010100",
    "1111001001110000",
    "1111011000101010",
    "1111101000001011",
    "1111111000101100",
    "1111110100010000",
    "1111011110101001",
    "1111001000100010",
    "1110110101000110",
    "1110101000001001",
    "1110100100101111",
    "1110101011001111",
    "1110111010100000",
    "1111010000100111",
    "1111101011010000",
    "1111110111100111",
    "1111011010000010",
    "1110111110011001",
    "1110100111001000",
    "1110010110101010",
    "1110001110110001",
    "1110001111100100",
    "1110011000011010",
    "1110101000110100",
    "1110111111110000",
    "1111011011011110",
    "1111111001010010",
    "1111101010001010",
    "1111010010010000",
    "1111000010000011",
    "1110111011011110",
    "1110111110001100",
    "1111000111100111",
    "1111010100000000",
    "1111100000010101",
    "1111101011111010",
    "1111110111110110",
    "1111111010100011",
    "1111101011001100",
    "1111011011111000",
    "1111010000001111",
    "1111001100100110",
    "1111010100100000",
    "1111101000111011",
    "1111111000101101",
    "1111010101100100",
    "1110110011100111",
    "1110011000001011",
    "1110000110100010",
    "1101111111100110",
    "1110000010001101",
    "1110001011111010",
    "1110011010011000",
    "1110101100010100",
    "1111000010000011",
    "1111011100011110",
    "1111111011110001",
    "1111100001011111",
    "1110111110010111",
    "1110011110001101",
    "1110000100010011",
    "1101110011001010",
    "1101101011110101",
    "1101101101100011",
    "1101110110001011",
    "1110000011000000",
    "1110010001011001",
    "1110011111000101",
    "1110101010101101",
    "1110110100011010",
    "1110111110001010",
    "1111001010010110",
    "1111011010000110",
    "1111101100011001",
    "1111111110011100",
    "1111110011001000",
    "1111101010110101",
    "1111101001001010",
    "1111101100000101",
    "1111101111110101",
    "1111110000101100",
    "1111101100100000",
    "1111100011100001",
    "1111010111110101",
    "1111001100001110",
    "1111000010101110",
    "1110111100010011",
    "1110111000101100",
    "1110110111001001",
    "1110110111000011",
    "1110111000010000",
    "1110111011000110",
    "1111000000010100",
    "1111001000000100",
    "1111010010001010",
    "1111011111111000",
    "1111110011100010",
    "1111110001101101",
    "1111010001001111",
    "1110101111001111",
    "1110010001010111",
    "1101111100101101",
    "1101110100011101",
    "1101111000011000",
    "1110000100011010",
    "1110010011000011",
    "1110011111011010",
    "1110100110111011",
    "1110101010000110",
    "1110101100111111",
    "1110110110000011",
    "1111001010001110",
    "1111101001111010",
    "1111101111011100",
    "1111001001101011",
    "1110101100100000",
    "1110011101000101",
    "1110011100001100",
    "1110100101011000",
    "1110110010011001",
    "1110111101111010",
    "1111000100111011",
    "1111000111010001",
    "1111000110011011",
    "1111000110101111",
    "1111001110100100",
    "1111100001111001",
    "1111111111101110",
    "1111011011000010",
    "1110110111100000",
    "1110011100001110",
    "1110001101111000",
    "1110001101001100",
    "1110010110001001",
    "1110100010101111",
    "1110101110001111",
    "1110110111111010",
    "1111000010110100",
    "1111010010010111",
    "1111100111111010",
    "1111111110001110",
    "1111100101001001",
    "1111010011101100",
    "1111010000001111",
    "1111011101101101",
    "1111111010000011",
    "1111100000110101",
    "1110111011000111",
    "1110011011111010",
    "1110000111011111",
    "1101111111101100",
    "1110000100001010",
    "1110010010001101",
    "1110100110000001",
    "1110111011111100",
    "1111010010110110",
    "1111101011111001",
    "1111110111110101",
    "1111011001000100",
    "1110111010101111",
    "1110100001000101",
    "1110010000010111",
    "1110001011110111",
    "1110010100001101",
    "1110100110100101",
    "1110111110000100",
    "1111010110011011",
    "1111101110111101",
    "1111110110011000",
    "1111010111111010",
    "1110110101111001",
    "1110010011101001",
    "1101110110101000",
    "1101100100101100",
    "1101100010000010",
    "1101101110110011",
    "1110000110111001",
    "1110100011111001",
    "1110111111011010",
    "1111010101100111",
    "1111100110000011",
    "1111110010011011",
    "1111111101101101",
    "1111110101011011",
    "1111100101111100",
    "1111010100111011",
    "1111000101000110",
    "1110111001101010",
    "1110110100101110",
    "1110110110010010",
    "1110111100100011",
    "1111000101001000",
    "1111001101101001",
    "1111010100000000",
    "1111010110011101",
    "1111010100001010",
    "1111001101010100",
    "1111000010110100",
    "1110110110001001",
    "1110101001010101",
    "1110011110100110",
    "1110010111110111",
    "1110010110001000",
    "1110011001010001",
    "1110100001011110",
    "1110110000000000",
    "1111000110100010",
    "1111100101011101",
    "1111110101010001",
    "1111001110010001",
    "1110101011011101",
    "1110010010101110",
    "1110000111111100",
    "1110001011010110",
    "1110011001010011",
    "1110101011111100",
    "1110111101100001",
    "1111001010101000",
    "1111010010100110",
    "1111010110100111",
    "1111011000111001",
    "1111011011011000",
    "1111011111011001",
    "1111100111001000",
    "1111110100111101",
    "1111110110010111",
    "1111011100001010",
    "1111000000001010",
    "1110100111111110",
    "1110011001110000",
    "1110011010111101",
    "1110101101000010",
    "1111001100001010",
    "1111110001011010",
    "1111101011000011",
    "1111001111110110",
    "1111000000011111",
    "1110111101010111",
    "1111000011110001",
    "1111001111001010",
    "1111011100101000",
    "1111101011110010",
    "1111111101100011",
    "1111101101010011",
    "1111010101110001",
    "1110111110101001",
    "1110101011110010",
    "1110100000011111",
    "1110011110000100",
    "1110100010101110",
    "1110101010110111",
    "1110110010011101",
    "1110110110110001",
    "1110110111011011",
    "1110110110111100",
    "1110111001011001",
    "1111000010101001",
    "1111010100001010",
    "1111101100000011",
    "1111111010001011",
    "1111100100001110",
    "1111010111000100",
    "1111010101001001",
    "1111011101101110",
    "1111101101111010",
    "1111111110000011",
    "1111101001010101",
    "1111010101011111",
    "1111000010101110",
    "1110110000111000",
    "1110100000001111",
    "1110010010001010",
    "1110001000110010",
    "1110000110010010",
    "1110001011111100",
    "1110011001010001",
    "1110101011111111",
    "1111000001000101",
    "1111010110101101",
    "1111101100101010",
    "1111111100011110",
    "1111100100100101",
    "1111001100101101",
    "1110110110111100",
    "1110100101111100",
    "1110011100000010",
    "1110011010011101",
    "1110100000101001",
    "1110101100111000",
    "1110111101000000",
    "1111001111010100",
    "1111100010111110",
    "1111110111101011",
    "1111110010110000",
    "1111011101001010",
    "1111001001000111",
    "1110111000100111",
    "1110101101001100",
    "1110100111100011",
    "1110100110110111",
    "1110101001001100",
    "1110101100100001",
    "1110101111010111",
    "1110110001001101",
    "1110110010010100",
    "1110110010111110",
    "1110110011011100",
    "1110110011101001",
    "1110110011011000",
    "1110110010110001",
    "1110110010001000",
    "1110110010000011",
    "1110110011001000",
    "1110110101010101",
    "1110111000000100",
    "1110111010011000",
    "1110111011100001",
    "1110111011110111",
    "1110111101110101",
    "1111000101111110",
    "1111011000000100",
    "1111110100110011",
    "1111100111010000",
    "1111000010101110",
    "1110100100100010",
    "1110010001111110",
    "1110001100110010",
    "1110010010001011",
    "1110011101000000",
    "1110101000010001",
    "1110110001011010",
    "1110111001100010",
    "1111000100000110",
    "1111010100011101",
    "1111101011111011",
    "1111110111010101",
    "1111011010001110",
    "1111000010001000",
    "1110110011010101",
    "1110101111011111",
    "1110110101010111",
    "1111000010011100",
    "1111010100100101",
    "1111101010100110",
    "1111111100001001",
    "1111100000111011",
    "1111000101101111",
    "1110101101001010",
    "1110011010000111",
    "1110001110111000",
    "1110001100000010",
    "1110010000011001",
    "1110011001001110",
    "1110100011001010",
    "1110101011001100",
    "1110101111110110",
    "1110110001001000",
    "1110110001000011",
    "1110110011100100",
    "1110111100001111",
    "1111001100001100",
    "1111100001001100",
    "1111110101111010",
    "1111111011111100",
    "1111111001101011",
    "1111111010010000",
    "1111100001111110",
    "1111000011100110",
    "1110100110111011",
    "1110010010111101",
    "1110001011100011",
    "1110010001010000",
    "1110100011011100",
    "1111000000101011",
    "1111100110011100",
    "1111101110101110",
    "1111000011110001",
    "1110011110001001",
    "1110000010011111",
    "1101110100000000",
    "1101110011001010",
    "1101111101010001",
    "1110001101110000",
    "1110011111101011",
    "1110101111100110",
    "1110111100011100",
    "1111000110101000",
    "1111001111011110",
    "1111011000001110",
    "1111100001011010",
    "1111101011111101",
    "1111111001110000",
    "1111110011101110",
    "1111011100011100",
    "1111000010010010",
    "1110101000111111",
    "1110010101001001",
    "1110001011000111",
    "1110001101001001",
    "1110011001101010",
    "1110101100010110",
    "1110111111111010",
    "1111001111110101",
    "1111011001100101",
    "1111011100111000",
    "1111011100000111",
    "1111011100101011",
    "1111100011110011",
    "1111110011101111",
    "1111110100111001",
    "1111011010110010",
    "1111000011010111",
    "1110110010110110",
    "1110101011010001",
    "1110101011010110",
    "1110101111101110",
    "1110110100111100",
    "1110111000110111",
    "1110111011000110",
    "1110111100101010",
    "1110111110100110",
    "1111000001100111",
    "1111000101110110",
    "1111001011100000",
    "1111010011111011",
    "1111100000010101",
    "1111110001000001",
    "1111111011010010",
    "1111100111011000",
    "1111010110101101",
    "1111001100011110",
    "1111001010000001",
    "1111001101100001",
    "1111010010111000",
    "1111010101111110",
    "1111010100010111",
    "1111001101110101",
    "1111000100000000",
    "1110111001011000",
    "1110110000101001",
    "1110101011110111",
    "1110101011100110",
    "1110101111001100",
    "1110110101011010",
    "1110111101000111",
    "1111000101111100",
    "1111010000000111",
    "1111011011111000",
    "1111101000111001",
    "1111110110010111",
    "1111111100110100",
    "1111110001100000",
    "1111101000001010",
    "1111100000111000",
    "1111011011011110",
    "1111010111111001",
    "1111010110010011",
    "1111010111001000",
    "1111011010110000",
    "1111100001010000",
    "1111101010001011",
    "1111110100101110",
    "1111111111110110",
    "1111110101101001",
    "1111101100111101",
    "1111100110110001",
    "1111100011000101",
    "1111100001100001",
    "1111100001100111",
    "1111100010110110",
    "1111100100100100",
    "1111100110000001",
    "1111100110100111",
    "1111100101111110",
    "1111100011111100",
    "1111100000100110",
    "1111011100100011",
    "1111011001000010",
    "1111010111100010",
    "1111011001011000",
    "1111011111010010",
    "1111101000111100",
    "1111110101001001",
    "1111111101101010",
    "1111110001000010",
    "1111100101110001",
    "1111011011110111",
    "1111010010110110",
    "1111001001111111",
    "1111000001001000",
    "1110111000100111",
    "1110110001011010",
    "1110101100101011",
    "1110101011000110",
    "1110101100111000",
    "1110110001100110",
    "1110111001011110",
    "1111000110010101",
    "1111011010011000",
    "1111110110010110",
    "1111100111011010",
    "1111000011010111",
    "1110100011010000",
    "1110001100100001",
    "1110000010100110",
    "1110000101001101",
    "1110010000101100",
    "1110100000001100",
    "1110101111001000",
    "1110111010111101",
    "1111000011010101",
    "1111001001000010",
    "1111001101100100",
    "1111010010000101",
    "1111010110101101",
    "1111011010101011",
    "1111011101000100",
    "1111011101010001",
    "1111011011101101",
    "1111011010000100",
    "1111011011001010",
    "1111100001110100",
    "1111101111011001",
    "1111111100101111",
    "1111100101100100",
    "1111001111001111",
    "1110111101111011",
    "1110110100101100",
    "1110110100010010",
    "1110111011001110",
    "1111000110111011",
    "1111010100111100",
    "1111100011100001",
    "1111110001100111",
    "1111111110011010",
    "1111110110110011",
    "1111101111000111",
    "1111101011100110",
    "1111101101001000",
    "1111110011101010",
    "1111111110010011",
    "1111110100011011",
    "1111100110011100",
    "1111011001011000",
    "1111001110011100",
    "1111000110001110",
    "1111000000111011",
    "1110111110110101",
    "1111000000111001",
    "1111001000101111",
    "1111010111110001",
    "1111101101110111",
    "1111110111001111",
    "1111011011100101",
    "1111000011100111",
    "1110110010111011",
    "1110101011011110",
    "1110101101001110",
    "1110110110110110",
    "1111000111000011",
    "1111011100111111",
    "1111110111111011",
    "1111101001110001",
    "1111001011001010",
    "1110110000001101",
    "1110011100110111",
    "1110010011101001",
    "1110010100110100",
    "1110011110001001",
    "1110101101000111",
    "1111000000110000",
    "1111011001010001",
    "1111110110110000",
    "1111101000011011",
    "1111001000000110",
    "1110101101001100",
    "1110011100101110",
    "1110011010000001",
    "1110100101001101",
    "1110111011011011",
    "1111011000010101",
    "1111110111100010",
    "1111101010001011",
    "1111001110101101",
    "1110110110110111",
    "1110100010111011",
    "1110010011010010",
    "1110001000101111",
    "1110000100001110",
    "1110000110111011",
    "1110010001110000",
    "1110100101001101",
    "1111000000011111",
    "1111100001011001",
    "1111111011101001",
    "1111011010110000",
    "1110111111110110",
    "1110101110000101",
    "1110100110110110",
    "1110101001011000",
    "1110110011001101",
    "1111000001001111",
    "1111010001001000",
    "1111100010001000",
    "1111110100001101",
    "1111111000110010",
    "1111100110001110",
    "1111010110100101",
    "1111001100111101",
    "1111001011111010",
    "1111010100010111",
    "1111100101000001",
    "1111111010101011",
    "1111101110100100",
    "1111011010000100",
    "1111001001100111",
    "1110111101100100",
    "1110110101100000",
    "1110110000101100",
    "1110101110101000",
    "1110101111010110",
    "1110110011010010",
    "1110111010111101",
    "1111000110110110",
    "1111010110111100",
    "1111101010110100",
    "1111111110101111",
    "1111101000000011",
    "1111010100001010",
    "1111000110100111",
    "1111000010101011",
    "1111001010010001",
    "1111011100111111",
    "1111110111101101",
    "1111101010010110",
    "1111001110100011",
    "1110111001001100",
    "1110101100110000",
    "1110101001110101",
    "1110110000001000",
    "1110111111001101",
    "1111010110011000",
    "1111110100000011",
    "1111101010100100",
    "1111001001011101",
    "1110101100110010",
    "1110011000001011",
    "1110001101100110",
    "1110001100111000",
    "1110010011111000",
    "1110011111101000",
    "1110101101110011",
    "1110111101001010",
    "1111001101011100",
    "1111011110100001",
    "1111101111110010",
    "1111111111110011",
    "1111110011001010",
    "1111101010101111",
    "1111100111001110",
    "1111100111011101",
    "1111101001010010",
    "1111101010011001",
    "1111101001011110",
    "1111100110101000",
    "1111100011000110",
    "1111100000011110",
    "1111011111110001",
    "1111100001001101",
    "1111100100010000",
    "1111101001010011",
    "1111110001111010",
    "1111111111100001",
    "1111101101101101",
    "1111010111110001",
    "1111000010010100",
    "1110110001100100",
    "1110101000111111",
    "1110101001100111",
    "1110110001000111",
    "1110111011001010",
    "1111000011100010",
    "1111000111011000",
    "1111000110110111",
    "1111000110000000",
    "1111001010110100",
    "1111011001100111",
    "1111110010100010",
    "1111101110110101",
    "1111010001100110",
    "1110111100010001",
    "1110110011001101",
    "1110110110100111",
    "1111000011010111",
    "1111010101111110",
    "1111101100000010",
    "1111111100001101",
    "1111100100011010",
    "1111001111000111",
    "1110111111011111",
    "1110111000010011",
    "1110111011110000",
    "1111001010011101",
    "1111100010100111",
    "1111111111001011",
    "1111011111111010",
    "1111000100100100",
    "1110110001001101",
    "1110101000000001",
    "1110101001010000",
    "1110110100000001",
    "1111000111000001",
    "1111100000010001",
    "1111111100111100",
    "1111100110010101",
    "1111001101000101",
    "1110111010000001",
    "1110101110010010",
    "1110101001100111",
    "1110101010110010",
    "1110110000110011",
    "1110111011000111",
    "1111001001100010",
    "1111011011100000",
    "1111101111111100",
    "1111111010100100",
    "1111100101100111",
    "1111010010011101",
    "1111000010010111",
    "1110110110101111",
    "1110110000111101",
    "1110110010010111",
    "1110111100000101",
    "1111001110011001",
    "1111101000001011",
    "1111111001001011",
    "1111011001101000",
    "1110111101100011",
    "1110101000111100",
    "1110011110011011",
    "1110011110111010",
    "1110101010001100",
    "1110111111001100",
    "1111011011110101",
    "1111111100110001",
    "1111100010010101",
    "1111000110001000",
    "1110110010010111",
    "1110101001000110",
    "1110101001111010",
    "1110110010011100",
    "1110111111100001",
    "1111001110110101",
    "1111011111101011",
    "1111110010101111",
    "1111110110111100",
    "1111011101011001",
    "1111000010001000",
    "1110101000100010",
    "1110010100110011",
    "1110001010001001",
    "1110001001101111",
    "1110010010001101",
    "1110100000010111",
    "1110110000101001",
    "1111000010000101",
    "1111010111010001",
    "1111110011011010",
    "1111101000101100",
    "1111000000000010",
    "1110011001000111",
    "1101111011011001",
    "1101101100110010",
    "1101101111011100",
    "1110000000000010",
    "1110010111101111",
    "1110110000110001",
    "1111001001000001",
    "1111100001011100",
    "1111111011100110",
    "1111101000111000",
    "1111001110101110",
    "1110111010001001",
    "1110101111110001",
    "1110110001100111",
    "1110111101100001",
    "1111001110000101",
    "1111011100111111",
    "1111100101011111",
    "1111100110011000",
    "1111100010001010",
    "1111011101110010",
    "1111011110110110",
    "1111101000101001",
    "1111111010110110",
    "1111101101111101",
    "1111010110111011",
    "1111000100110100",
    "1110111010100011",
    "1110111000010101",
    "1110111100000111",
    "1111000011000110",
    "1111001010110010",
    "1111010001110001",
    "1111011000110000",
    "1111100001101110",
    "1111101110101000",
    "1111111111111001",
    "1111101100011101",
    "1111011010011000",
    "1111001101111101",
    "1111001010001001",
    "1111001111110110",
    "1111011101011001",
    "1111101111110011",
    "1111111011111100",
    "1111100111111100",
    "1111010100111110",
    "1111000011100010",
    "1110110100001110",
    "1110100111110100",
    "1110011111001111",
    "1110011011100001",
    "1110011101101011",
    "1110100110101100",
    "1110110111010011",
    "1111001111011110",
    "1111101110000000",
    "1111101111101100",
    "1111001101011100",
    "1110101111011001",
    "1110011001100010",
    "1110001110101001",
    "1110001111011001",
    "1110011010000001",
    "1110101011011101",
    "1111000001000111",
    "1111011001111111",
    "1111110101110000",
    "1111101100010001",
    "1111001110001010",
    "1110110011100110",
    "1110100001000101",
    "1110011010110000",
    "1110100010101011",
    "1110110111010011",
    "1111010011110001",
    "1111110001010111",
    "1111110110101110",
    "1111101001101010",
    "1111101001100100",
    "1111110101001110",
    "1111110111000101",
    "1111100000010111",
    "1111001010111111",
    "1110111001111010",
    "1110101110001111",
    "1110100111011010",
    "1110100100000001",
    "1110100010101001",
    "1110100010010111",
    "1110100100011101",
    "1110101100100110",
    "1110111110010010",
    "1111011010101000",
    "1111111110111101",
    "1111011010100110",
    "1110111000110101",
    "1110100001001101",
    "1110010110000001",
    "1110010101010101",
    "1110011010110000",
    "1110100001101100",
    "1110100111011000",
    "1110101011011101",
    "1110101111001010",
    "1110110011111001",
    "1110111010111000",
    "1111000101000101",
    "1111010011011010",
    "1111100110011110",
    "1111111101011111",
    "1111101001111000",
    "1111010011010000",
    "1111000010100110",
    "1110111011001110",
    "1110111110100110",
    "1111001011000001",
    "1111011011111101",
    "1111101011111000",
    "1111110110011000",
    "1111111001101101",
    "1111110110101100",
    "1111101111100100",
    "1111100110100101",
    "1111011100110010",
    "1111010001111011",
    "1111000101011000",
    "1110110111001101",
    "1110101000110100",
    "1110011100110010",
    "1110010101111100",
    "1110010101111100",
    "1110011100010100",
    "1110100110111100",
    "1110110010111101",
    "1110111101111000",
    "1111000110101111",
    "1111001111111011",
    "1111011110100011",
    "1111110110011110",
    "1111101000000111",
    "1111000001101011",
    "1110011101110101",
    "1110000100001011",
    "1101111001111001",
    "1101111111110000",
    "1110010001010101",
    "1110100111101100",
    "1110111100011001",
    "1111001011011110",
    "1111010100100100",
    "1111011001110101",
    "1111011110011011",
    "1111100101010010",
    "1111101111011100",
    "1111111011111010",
    "1111110111010100",
    "1111101100100010",
    "1111100100111110",
    "1111100000001100",
    "1111011100101101",
    "1111011001000110",
    "1111010100110111",
    "1111010000101011",
    "1111001101101000",
    "1111001101000010",
    "1111010000000000",
    "1111010111011010",
    "1111100011100100",
    "1111110100010111",
    "1111110111000011",
    "1111100000100001",
    "1111001010011011",
    "1110110111101111",
    "1110101011000111",
    "1110100110000110",
    "1110101000101000",
    "1110110001000011",
    "1110111100101011",
    "1111001000111010",
    "1111010100100101",
    "1111100000010111",
    "1111101101111101",
    "1111111110010100",
    "1111101111010010",
    "1111011101011110",
    "1111001111001111",
    "1111000110110001",
    "1111000100011010",
    "1111000110100100",
    "1111001010100101",
    "1111001110000100",
    "1111001111101110",
    "1111001111101011",
    "1111001110110110",
    "1111001110011011",
    "1111001110111010",
    "1111001111110001",
    "1111010000000000",
    "1111001110100100",
    "1111001011010011",
    "1111000110110100",
    "1111000010101001",
    "1111000000100001",
    "1111000001101100",
    "1111000110110111",
    "1111010001011111",
    "1111100011011000",
    "1111111101010010",
    "1111100010001010",
    "1110111110111000",
    "1110011101111101",
    "1110000100000110",
    "1101110100110001",
    "1101110000101110",
    "1101110101101010",
    "1101111111111010",
    "1110001100001001",
    "1110011000011011",
    "1110100100100101",
    "1110110001001100",
    "1110111110110000",
    "1111001101101000",
    "1111011101001100",
    "1111101100001010",
    "1111111001010111",
    "1111111011111010",
    "1111110011100111",
    "1111101100110110",
    "1111100110100110",
    "1111100000011100",
    "1111011010110000",
    "1111010110000001",
    "1111010010011111",
    "1111010000001010",
    "1111001111000000",
    "1111001111001000",
    "1111010000100111",
    "1111010011101111",
    "1111011000111111",
    "1111100000111011",
    "1111101011110000",
    "1111111000101111",
    "1111111001101101",
    "1111101101101110",
    "1111100101001011",
    "1111100001000101",
    "1111100001011100",
    "1111100101010000",
    "1111101010110101",
    "1111110000100100",
    "1111110101010011",
    "1111111000010101",
    "1111111001000101",
    "1111110110110010",
    "1111110000110111",
    "1111100111100111",
    "1111011100100001",
    "1111010010010100",
    "1111001100001111",
    "1111001101011100",
    "1111010111110100",
    "1111101011001001",
    "1111111011000010",
    "1111011111000000",
    "1111000101011010",
    "1110110010000011",
    "1110100111001000",
    "1110100100111110",
    "1110101010001100",
    "1110110100010101",
    "1111000000101110",
    "1111001101001111",
    "1111011001110010",
    "1111101000110010",
    "1111111101001111",
    "1111100111011010",
    "1111000110100010",
    "1110100100001000",
    "1110000101011000",
    "1101101111000111",
    "1101100100010000",
    "1101100100001101",
    "1101101011011110",
    "1101110101101110",
    "1101111111010100",
    "1110000110011011",
    "1110001010111111",
    "1110001101111011",
    "1110010000111000",
    "1110010101000101",
    "1110011010110111",
    "1110100001110011",
    "1110101001011101",
    "1110110011100010",
    "1111000011110001",
    "1111011100101000",
    "1111111101100100",
    "1111011101101001",
    "1110111011101111",
    "1110100010101110",
    "1110010110100100",
    "1110010111101100",
    "1110100010110001",
    "1110110011001101",
    "1111000101010111",
    "1111010111001011",
    "1111101000011001",
    "1111111000111111",
    "1111110111101011",
    "1111101010100100",
    "1111100001000010",
    "1111011100000111",
    "1111011011100110",
    "1111011110011011",
    "1111100011000011",
    "1111100111111100",
    "1111101100001011",
    "1111101111101100",
    "1111110010101101",
    "1111110100111001",
    "1111110100111011",
    "1111110001010011",
    "1111101001011110",
    "1111011110011100",
    "1111010010011101",
    "1111001000011110",
    "1111000010111101",
    "1111000011001011",
    "1111001001100011",
    "1111010101101110",
    "1111100111000000",
    "1111111100011100",
    "1111101011000000",
    "1111010000101011",
    "1110110110100101",
    "1110011111010110",
    "1110001101100001",
    "1110000010111001",
    "1101111111110011",
    "1110000011000110",
    "1110001010101101",
    "1110010100000110",
    "1110011101110111",
    "1110101000110000",
    "1110110111001001",
    "1111001010111000",
    "1111100100000000",
    "1111111111110011",
    "1111100101110110",
    "1111010001001100",
    "1111000100101111",
    "1111000000010001",
    "1111000000110001",
    "1111000010000101",
    "1111000000100110",
    "1110111010111101",
    "1110110010010010",
    "1110101001010000",
    "1110100010111001",
    "1110100001011010",
    "1110100101010010",
    "1110101101100000",
    "1110110111111100",
    "1111000010010000",
    "1111001010110010",
    "1111010001000000",
    "1111010101011000",
    "1111011001001100",
    "1111011110010001",
    "1111100110011110",
    "1111110011100000",
    "1111111010000000",
    "1111100011010111",
    "1111001011000100",
    "1110110100010010",
    "1110100001101100",
    "1110010100101111",
    "1110001101011001",
    "1110001010010100",
    "1110001001101000",
    "1110001001110100",
    "1110001010011101",
    "1110001100001100",
    "1110010000100100",
    "1110011001111100",
    "1110101011000010",
    "1111000101011010",
    "1111101000000101",
    "1111110000111010",
    "1111001011101000",
    "1110101110001001",
    "1110011100110101",
    "1110011001001011",
    "1110100001000101",
    "1110110000000010",
    "1111000000101011",
    "1111001110101000",
    "1111011000000100",
    "1111011111011100",
    "1111101001011110",
    "1111111001111110",
    "1111101110011101",
    "1111010011101001",
    "1110111011111111",
    "1110101110000101",
    "1110101110101011",
    "1110111110000101",
    "1111010111100010",
    "1111110100000010",
    "1111110011001001",
    "1111100010010000",
    "1111011010000111",
    "1111011001011110",
    "1111011101101000",
    "1111100011100111",
    "1111101010000011",
    "1111110001001111",
    "1111111010011111",
    "1111111000110111",
    "1111101000101111",
    "1111010110101010",
    "1111000100111011",
    "1110110101100010",
    "1110101001111111",
    "1110100011000101",
    "1110100001001100",
    "1110100011110110",
    "1110101001110101",
    "1110110001011111",
    "1110111001001110",
    "1110111111101100",
    "1111000100000000",
    "1111000110101000",
    "1111001010110101",
    "1111010101000101",
    "1111100111100101",
    "1111111110111100",
    "1111100011101010",
    "1111001101011100",
    "1111000010010000",
    "1111000101011111",
    "1111010101111001",
    "1111101101110010",
    "1111111010000110",
    "1111100111110101",
    "1111011110001010",
    "1111011100000100",
    "1111011100111010",
    "1111011001110101",
    "1111001101101101",
    "1110110111111111",
    "1110011100110010",
    "1110000010111110",
    "1101110001011110",
    "1101101100111000",
    "1101110101100101",
    "1110000111011000",
    "1110011101000111",
    "1110110100010000",
    "1111001100101000",
    "1111100111000100",
    "1111111100011110",
    "1111100000010001",
    "1111000111110100",
    "1110110111100111",
    "1110110011101100",
    "1110111101000111",
    "1111010001100010",
    "1111101100001010",
    "1111111000111011",
    "1111100010110110",
    "1111010100101111",
    "1111001111110001",
    "1111010011011010",
    "1111011110001111",
    "1111101110010000",
    "1111111111010000",
    "1111101101110001",
    "1111100000101110",
    "1111011011000110",
    "1111011110100100",
    "1111101010110101",
    "1111111101011000",
    "1111101101011101",
    "1111011001110000",
    "1111001010101011",
    "1111000010001010",
    "1111000000101001",
    "1111000100101010",
    "1111001011011001",
    "1111010001100001",
    "1111010100011000",
    "1111010011000101",
    "1111001110000000",
    "1111000110111001",
    "1111000000000000",
    "1110111011100011",
    "1110111011000010",
    "1110111111001101",
    "1111001000101100",
    "1111011000010011",
    "1111101110001000",
    "1111110111010111",
    "1111011011100001",
    "1111000010100111",
    "1110110000100001",
    "1110100111100111",
    "1110100111111100",
    "1110101111001010",
    "1110111010001001",
    "1111000110110100",
    "1111010100111110",
    "1111100101101111",
    "1111111010000010",
    "1111101110111111",
    "1111011000001011",
    "1111000101010101",
    "1110111001111100",
    "1110110111011011",
    "1110111100111000",
    "1111001000001001",
    "1111010110111001",
    "1111100111100011",
    "1111111001011101",
    "1111110100000100",
    "1111100010101111",
    "1111010101100111",
    "1111010000011110",
    "1111010110010011",
    "1111100111011110",
    "1111111111000111",
    "1111100011001101",
    "1111001011000010",
    "1110111011100001",
    "1110110110100101",
    "1110111011000111",
    "1111000101110010",
    "1111010011001000",
    "1111100011000110",
    "1111111000100110",
    "1111101010000001",
    "1111000101000011",
    "1110011100100110",
    "1101110111101010",
    "1101011101000101",
    "1101010001100110",
    "1101010101011010",
    "1101100011101010",
    "1101110101100010",
    "1110000101000110",
    "1110001111000101",
    "1110010011101100",
    "1110010100110111",
    "1110010100101111",
    "1110010101001001",
    "1110010110100000",
    "1110011000100101",
    "1110011100100011",
    "1110100100111011",
    "1110110100000011",
    "1111001010100110",
    "1111100101111110",
    "1111111111011100",
    "1111101100001100",
    "1111100101001000",
    "1111101011001110",
    "1111111011000110",
    "1111110000111011",
    "1111011110110011",
    "1111010010101110",
    "1111001101111101",
    "1111001111101100",
    "1111010101111001",
    "1111011110010010",
    "1111100111011010",
    "1111110000110110",
    "1111111010011100",
    "1111111011110111",
    "1111110010011110",
    "1111101010000001",
    "1111100011000011",
    "1111011101101000",
    "1111011001001001",
    "1111010100110111",
    "1111010000101011",
    "1111001101001110",
    "1111001011100000",
    "1111001100100001",
    "1111010000110101",
    "1111011000011101",
    "1111100011001000",
    "1111110000000100",
    "1111111101110111",
    "1111110101010010",
    "1111101011101000",
    "1111100111000111",
    "1111101001000101",
    "1111110001110011",
    "1111111111101001",
    "1111101101100110",
    "1111011011000010",
    "1111001011010100",
    "1111000001010100",
    "1110111110110110",
    "1111000100110011",
    "1111010011010000",
    "1111101001101011",
    "1111111001011000",
    "1111011000100010",
    "1110110111010110",
    "1110011010000110",
    "1110000100100100",
    "1101111000110111",
    "1101110110100010",
    "1101111010110000",
    "1110000001110000",
    "1110001000000100",
    "1110001100101010",
    "1110010001011100",
    "1110011010001111",
    "1110101010001111",
    "1111000010011001",
    "1111100000010100",
    "1111111111001100",
    "1111100110010110",
    "1111010100100111",
    "1111001100110011",
    "1111001101001111",
    "1111010010101011",
    "1111011001101101",
    "1111100000001101",
    "1111100101001110",
    "1111101000101010",
    "1111101010101100",
    "1111101011001111",
    "1111101001101011",
    "1111100101001110",
    "1111011101100001",
    "1111010010111110",
    "1111000111000001",
    "1110111011101101",
    "1110110010111101",
    "1110101101110101",
    "1110101100011011",
    "1110101110001100",
    "1110110010011001",
    "1110111000011010",
    "1110111111110101",
    "1111001000100010",
    "1111010010110001",
    "1111011111011001",
    "1111101111110011",
    "1111111010110111",
    "1111100000110001",
    "1111000011110100",
    "1110100111101000",
    "1110010000101001",
    "1110000010101100",
    "1101111111101110",
    "1110000110110110",
    "1110010100110110",
    "1110100101011010",
    "1110110100011000",
    "1110111111110000",
    "1111001001101010",
    "1111010110111001",
    "1111101011000110",
    "1111111001011000",
    "1111011010101010",
    "1110111111100110",
    "1110101111010001",
    "1110101111001000",
    "1111000000010111",
    "1111011110111010",
    "1111111100000011",
    "1111011000001000",
    "1110111011010110",
    "1110101000111010",
    "1110100001110000",
    "1110100100100100",
    "1110101110101110",
    "1110111101101011",
    "1111001111001100",
    "1111100001001100",
    "1111110001100111",
    "1111111110001001",
    "1111111011100011",
    "1111111100111000",
    "1111111010101110",
    "1111101101111000",
    "1111100000010100",
    "1111010101110111",
    "1111010010000010",
    "1111010111000100",
    "1111100101010000",
    "1111111010011010",
    "1111101101001010",
    "1111010110001000",
    "1111000100010011",
    "1110111001110100",
    "1110110110101111",
    "1110111001011000",
    "1110111110111101",
    "1111000100101100",
    "1111001000100011",
    "1111001001110100",
    "1111001001010110",
    "1111001001101010",
    "1111001101101101",
    "1111010111011111",
    "1111100110100110",
    "1111111000100101",
    "1111110110001010",
    "1111101001000100",
    "1111100010000101",
    "1111100001010101",
    "1111100101100100",
    "1111101101010111",
    "1111110111101010",
    "1111111100001100",
    "1111101110111011",
    "1111100001100111",
    "1111010101110110",
    "1111001101110101",
    "1111001100000111",
    "1111010010011101",
    "1111100001001010",
    "1111110110011011",
    "1111110001001100",
    "1111011010000010",
    "1111000111111010",
    "1110111101001111",
    "1110111010100110",
    "1110111111001100",
    "1111001001010011",
    "1111010111000110",
    "1111100110101110",
    "1111110110010010",
    "1111111100000101",
    "1111110010001001",
    "1111101101001101",
    "1111101101100011",
    "1111110010001111",
    "1111111001000000",
    "1111111110101111",
    "1111111111011001",
    "1111111100110011",
    "1111110011101010",
    "1111100111001000",
    "1111011010000110",
    "1111001111010111",
    "1111001000110101",
    "1111000110111100",
    "1111001000111100",
    "1111001101011100",
    "1111010010111110",
    "1111011000011110",
    "1111011101011001",
    "1111100001110100",
    "1111100110011000",
    "1111101011101110",
    "1111110010001101",
    "1111111001110011",
    "1111111101111011",
    "1111110101100110",
    "1111101101100000",
    "1111100101110110",
    "1111011110101110",
    "1111011000010101",
    "1111010011001011",
    "1111001111111011",
    "1111001111010100",
    "1111010001111000",
    "1111010111101101",
    "1111100000011010",
    "1111101011001111",
    "1111110111011001",
    "1111111011111101",
    "1111101111111001",
    "1111100101011000",
    "1111011101100000",
    "1111011000111111",
    "1111011000001110",
    "1111011011000010",
    "1111100000101100",
    "1111101000001100",
    "1111110000111011",
    "1111111010111101",
    "1111111001011001",
    "1111101100011000",
    "1111011111001100",
    "1111010100000000",
    "1111001101101011",
    "1111001110111111",
    "1111011010001001",
    "1111101111110011",
    "1111110001100000",
    "1111001101100000",
    "1110101001001100",
    "1110001010000110",
    "1101110100100000",
    "1101101010110010",
    "1101101100101010",
    "1101110111010110",
    "1110000111010101",
    "1110011010111010",
    "1110110010111110",
    "1111010000111000",
    "1111110100011011",
    "1111100101011010",
    "1111000001111110",
    "1110100110111011",
    "1110011000101111",
    "1110011000101101",
    "1110100011111000",
    "1110110100101100",
    "1111000101011111",
    "1111010010001111",
    "1111011001110010",
    "1111011100111000",
    "1111011101000111",
    "1111011100001111",
    "1111011011001010",
    "1111011010000110",
    "1111011001101101",
    "1111011011110111",
    "1111100011100110",
    "1111110011010100",
    "1111110100110000",
    "1111010111101111",
    "1110111010110101",
    "1110100011101110",
    "1110010110001001",
    "1110010010110011",
    "1110010111010000",
    "1110011111010001",
    "1110100110111111",
    "1110101101101001",
    "1110110101101111",
    "1111000010011111",
    "1111010101110001",
    "1111101110001111",
    "1111111000011000",
    "1111100011100010",
    "1111010111101111",
    "1111010110100000",
    "1111011101010001",
    "1111100111000101",
    "1111101110111011",
    "1111110001110101",
    "1111110000000110",
    "1111101100101000",
    "1111101011111001",
    "1111110001101000",
    "1111111110100001",
    "1111110000010001",
    "1111100000010001",
    "1111010111011010",
    "1111011010000100",
    "1111101001010110",
    "1111111101110000",
    "1111100001000000",
    "1111000110101000",
    "1110110011100111",
    "1110101010111010",
    "1110101110000010",
    "1110111101011110",
    "1111011000000110",
    "1111111010111001",
    "1111011110100001",
    "1110111001101010",
    "1110011011101011",
    "1110001000010110",
    "1110000001000011",
    "1110000100000000",
    "1110001101001001",
    "1110010111110001",
    "1110100000010111",
    "1110100101101010",
    "1110101000100000",
    "1110101010111101",
    "1110101111011001",
    "1110111000011010",
    "1111000111110010",
    "1111011101111111",
    "1111111001110000",
    "1111100111111011",
    "1111001011001010",
    "1110110011111011",
    "1110100101011111",
    "1110100001000101",
    "1110100101101111",
    "1110110001000000",
    "1110111111101110",
    "1111001111000100",
    "1111011100110101",
    "1111100111011011",
    "1111101101111110",
    "1111110000011101",
    "1111101111011001",
    "1111101011111011",
    "1111100111110101",
    "1111100101001011",
    "1111100110001101",
    "1111101100011000",
    "1111110111110110",
    "1111111000110011",
    "1111101000011001",
    "1111011001101111",
    "1111001110101101",
    "1111000111101111",
    "1111000011111110",
    "1111000010000011",
    "1111000000110001",
    "1110111111011001",
    "1110111101101101",
    "1110111011111101",
    "1110111010110100",
    "1110111010101101",
    "1110111011110111",
    "1110111110010001",
    "1111000001111101",
    "1111000111111100",
    "1111010010010000",
    "1111100010010100",
    "1111110111101111",
    "1111110000100101",
    "1111011100010110",
    "1111010001111110",
    "1111010110011011",
    "1111101010110110",
    "1111110100101111",
    "1111010000000111",
    "1110101111110000",
    "1110011010010011",
    "1110010010100001",
    "1110010111010011",
    "1110100100101010",
    "1110110101010011",
    "1111000100110011",
    "1111010000101011",
    "1111011001011001",
    "1111100010001101",
    "1111101110101101",
    "1111111111100011",
    "1111101001111110",
    "1111010100010010",
    "1111000010100111",
    "1110111000001100",
    "1110110110010110",
    "1110111011011001",
    "1111000011011111",
    "1111001010011011",
    "1111001101001001",
    "1111001010110000",
    "1111000100011111",
    "1110111100100101",
    "1110110110010000",
    "1110110100111100",
    "1110111010111111",
    "1111001000111110",
    "1111011101000100",
    "1111110011011011",
    "1111111000011101",
    "1111101010011011",
    "1111100100011100",
    "1111100110000000",
    "1111101100011000",
    "1111110011100110",
    "1111111000011000",
    "1111111010100001",
    "1111111100111001",
    "1111111100111101",
    "1111110001010010",
    "1111100001011110",
    "1111010001111001",
    "1111001000001001",
    "1111001000111010",
    "1111010110010101",
    "1111101110100010",
    "1111110011001110",
    "1111010101000001",
    "1110111011111000",
    "1110101010100110",
    "1110100010000010",
    "1110100001100001",
    "1110100111011111",
    "1110110010000110",
    "1111000000000000",
    "1111010000111000",
    "1111100101110111",
    "1111111111101101",
    "1111100000000111",
    "1110111101001111",
    "1110011010011011",
    "1101111011100001",
    "1101100100000000",
    "1101010110011000",
    "1101010011001101",
    "1101011001011001",
    "1101101000000001",
    "1101111110110101",
    "1110011101010100",
    "1111000001100110",
    "1111100111100100",
    "1111110110011010",
    "1111011101110011",
    "1111010010111000",
    "1111010111010000",
    "1111101001010000",
    "1111111011010001",
    "1111011011111101",
    "1110111110001100",
    "1110100101110110",
    "1110010101110010",
    "1110010000000101",
    "1110010110000001",
    "1110100111100111",
    "1111000010110001",
    "1111100011000110",
    "1111111100110100",
    "1111100010011101",
    "1111010001101110",
    "1111001011101010",
    "1111001110010100",
    "1111010101011111",
    "1111011100111100",
    "1111100001111000",
    "1111100011111110",
    "1111100110010011",
    "1111101110010100",
    "1111111111011001",
    "1111100001101001",
    "1110111011101000",
    "1110010100000101",
    "1101110010110011",
    "1101011110001100",
    "1101011000111010",
    "1101100001000000",
    "1101110001110100",
    "1110000110100010",
    "1110011011010100",
    "1110101110010100",
    "1110111110110000",
    "1111001100010110",
    "1111011000001100",
    "1111100100111100",
    "1111110100110100",
    "1111110111011101",
    "1111100001011110",
    "1111001101000000",
    "1110111110010111",
    "1110111001011011",
    "1111000000101100",
    "1111010100000000",
    "1111110000010010",
    "1111101111011000",
    "1111010001000000",
    "1110111001100000",
    "1110101011101011",
    "1110101000001011",
    "1110101100111101",
    "1110110110100010",
    "1111000010110100",
    "1111010010011100",
    "1111100110110010",
    "1111111111101001",
    "1111100011001101",
    "1111001000101010",
    "1110110101010111",
    "1110101101100011",
    "1110110010111101",
    "1111000011110001",
    "1111011100111101",
    "1111111011100000",
    "1111100011101110",
    "1111000011110001",
    "1110100111111111",
    "1110010100000110",
    "1110001010111101",
    "1110001110110001",
    "1110100000000111",
    "1110111100101101",
    "1111100000001100",
    "1111111010110101",
    "1111011001110010",
    "1111000000011010",
    "1110110000011111",
    "1110101001000001",
    "1110100110111111",
    "1110100111001000",
    "1110100110111110",
    "1110100101010011",
    "1110100010010100",
    "1110011111001100",
    "1110011101101000",
    "1110011111000010",
    "1110100100010010",
    "1110101100111010",
    "1110110111010101",
    "1111000001011110",
    "1111001001100011",
    "1111001111011001",
    "1111010110001001",
    "1111100010100111",
    "1111110111110001",
    "1111101010111010",
    "1111001010000100",
    "1110101100011110",
    "1110011000011101",
    "1110010010001111",
    "1110011001101010",
    "1110101010000100",
    "1110111101000100",
    "1111001100101101",
    "1111010101100111",
    "1111010111110100",
    "1111010101011111",
    "1111010001110100",
    "1111001111110101",
    "1111010000110001",
    "1111010100100000",
    "1111011011000001",
    "1111100100100100",
    "1111110001111100",
    "1111111100000001",
    "1111100101111001",
    "1111001101111101",
    "1110110111101101",
    "1110100110100111",
    "1110011100010100",
    "1110011000001001",
    "1110010111111111",
    "1110011001001011",
    "1110011001101010",
    "1110011001000010",
    "1110011000001001",
    "1110011000100101",
    "1110011100101010",
    "1110100110111100",
    "1110111001101000",
    "1111010101001001",
    "1111110111011111",
    "1111100011100111",
    "1111000001110000",
    "1110101000000100",
    "1110011010000010",
    "1110011000000100",
    "1110011111011110",
    "1110101011100110",
    "1110110111011010",
    "1110111111100001",
    "1111000100010111",
    "1111001001100000",
    "1111010011000011",
    "1111100011010000",
    "1111111001000000",
    "1111101111110111",
    "1111011100110000",
    "1111010010010000",
    "1111010010010100",
    "1111011011001111",
    "1111101001000100",
    "1111110111001110",
    "1111111101100111",
    "1111110110101110",
    "1111110011110011",
    "1111110011110010",
    "1111110101011010",
    "1111111000010111",
    "1111111101100110",
    "1111111001011111",
    "1111101011111110",
    "1111011010000111",
    "1111000101110010",
    "1110110001110000",
    "1110100000100100",
    "1110010100010101",
    "1110001101111101",
    "1110001101100100",
    "1110010010101001",
    "1110011100001111",
    "1110101001000110",
    "1110111000000011",
    "1111001000001001",
    "1111011001010101",
    "1111101100001001",
    "1111111111000101",
    "1111101001000011",
    "1111010011110100",
    "1111000010100010",
    "1110111000010000",
    "1110110110111011",
    "1110111110011100",
    "1111001100110000",
    "1111011111100001",
    "1111110110000101",
    "1111101110111101",
    "1111001111011111",
    "1110101100111010",
    "1110001011000001",
    "1101101111000100",
    "1101011110001100",
    "1101011011100101",
    "1101100110011111",
    "1101111010000111",
    "1110010000010100",
    "1110100011011000",
    "1110110000110001",
    "1110111010111010",
    "1111000111010011",
    "1111011010111111",
    "1111110111111011",
    "1111100100110100",
    "1111000001100110",
    "1110100101001000",
    "1110010100110100",
    "1110010001101100",
    "1110011000001100",
    "1110100010111000",
    "1110101100111100",
    "1110110011110100",
    "1110110111010110",
    "1110111000010110",
    "1110111000001000",
    "1110111000001001",
    "1110111000111001",
    "1110111010010011",
    "1110111101100000",
    "1111000101010010",
    "1111010100011111",
    "1111101100001010",
    "1111110101110101",
    "1111010110100111",
    "1110111100000001",
    "1110101010101011",
    "1110100100010111",
    "1110100110111111",
    "1110101110011011",
    "1110110110100111",
    "1110111100111111",
    "1111000000111110",
    "1111000010111011",
    "1111000011000101",
    "1111000001100110",
    "1110111110011100",
    "1110111001101010",
    "1110110100000011",
    "1110101111000101",
    "1110101100010011",
    "1110101101000000",
    "1110110001101100",
    "1110111001110100",
    "1111000011111011",
    "1111001111001010",
    "1111011100011011",
    "1111101101100110",
    "1111111100010011",
    "1111100010101110",
    "1111001001001100",
    "1110110100001011",
    "1110100111100000",
    "1110100100111011",
    "1110101011110010",
    "1110111001110111",
    "1111001100110011",
    "1111100010110110",
    "1111111010110101",
    "1111101100010110",
    "1111010100001101",
    "1110111110100001",
    "1110101101100000",
    "1110100011000011",
    "1110100000000011",
    "1110100011111001",
    "1110101100101110",
    "1110111000011101",
    "1111000101100100",
    "1111010011111011",
    "1111100100010101",
    "1111110111010111",
    "1111110011110010",
    "1111011111101001",
    "1111001111010110",
    "1111000101001110",
    "1111000001111110",
    "1111000100001000",
    "1111001000111001",
    "1111001101000000",
    "1111001101111010",
    "1111001010010100",
    "1111000010010010",
    "1110110110101111",
    "1110101001010110",
    "1110011100001001",
    "1110010001000101",
    "1110001001101010",
    "1110000110011111",
    "1110000111001011",
    "1110001010101111",
    "1110001111101011",
    "1110010100100010",
    "1110011000010101",
    "1110011011001010",
    "1110011110010100",
    "1110100011011000",
    "1110101011101010",
    "1110110111010000",
    "1111000100111100",
    "1111010010101001",
    "1111011110001100",
    "1111100110011001",
    "1111101011011010",
    "1111101110111100",
    "1111110011100000",
    "1111111011001000",
    "1111111001101111",
    "1111101100111000",
    "1111100001010010",
    "1111011001111100",
    "1111011000101000",
    "1111011101001111",
    "1111100101110010",
    "1111101111011111",
    "1111110111110101",
    "1111111110000010",
    "1111111101000111",
    "1111111000011111",
    "1111110011100011",
    "1111101111001111",
    "1111101101110001",
    "1111110001011011",
    "1111111011011101",
    "1111110100101110",
    "1111100010000101",
    "1111010000100011",
    "1111000011100100",
    "1110111100101101",
    "1110111011101011",
    "1110111111111000",
    "1111001001000110",
    "1111010111001101",
    "1111101001011101",
    "1111111101111001",
    "1111101110010110",
    "1111011110101011",
    "1111010101101110",
    "1111010100100100",
    "1111011010001001",
    "1111100011110100",
    "1111101110011110",
    "1111110111011010",
    "1111111101000000",
    "1111111110100000",
    "1111111011101011",
    "1111110100111000",
    "1111101010110000",
    "1111011110010111",
    "1111010001010010",
    "1111000101110100",
    "1110111111000000",
    "1111000000000101",
    "1111001010110010",
    "1111011110001100",
    "1111110110011011",
    "1111110010000011",
    "1111100000100001",
    "1111011000001100",
    "1111011001100101",
    "1111100010011001",
    "1111101110110101",
    "1111111011001011",
    "1111111011001000",
    "1111110101000111",
    "1111110010110001",
    "1111110011111010",
    "1111111000101100",
    "1111111110001101",
    "1111110000001100",
    "1111011101100001",
    "1111000111110001",
    "1110110001011110",
    "1110011101111010",
    "1110001111111010",
    "1110001000111110",
    "1110001000110101",
    "1110001101111000",
    "1110010101110001",
    "1110011110011011",
    "1110100110010110",
    "1110101100110111",
    "1110110001111011",
    "1110110110001000",
    "1110111010010100",
    "1111000000010001",
    "1111001010011101",
    "1111011010111101",
    "1111110010001001",
    "1111110010000111",
    "1111010110010000",
    "1110111111001000",
    "1110110000100110",
    "1110101100000100",
    "1110101111110000",
    "1110110111100010",
    "1110111110110001",
    "1111000001111000",
    "1110111111010111",
    "1110111000000100",
    "1110101110001010",
    "1110100100011111",
    "1110011101010010",
    "1110011001101010",
    "1110011001100101",
    "1110011100100001",
    "1110100001111101",
    "1110101010000001",
    "1110110101100100",
    "1111000100111001",
    "1111010111010001",
    "1111101010100110",
    "1111111100010110",
    "1111110101011011",
    "1111101011101110",
    "1111100110000000",
    "1111100010011101",
    "1111011110101101",
    "1111011000100011",
    "1111001111000010",
    "1111000010101111",
    "1110110101100010",
    "1110101001110010",
    "1110100001111110",
    "1110100000010101",
    "1110100110101010",
    "1110110101110110",
    "1111001101000111",
    "1111101001111111",
    "1111110111100010",
    "1111011100001110",
    "1111001000001001",
    "1110111101101101",
    "1110111100110010",
    "1111000011000000",
    "1111001100110011",
    "1111010110110110",
    "1111011110110001",
    "1111100100010000",
    "1111101001010101",
    "1111110001001000",
    "1111111101111100",
    "1111110000010011",
    "1111011100100001",
    "1111001010111111",
    "1110111111111011",
    "1110111110010111",
    "1111000111001101",
    "1111011001001011",
    "1111110001100110",
    "1111110011000000",
    "1111011000010000",
    "1111000001010101",
    "1110110001001000",
    "1110101010011011",
    "1110101111111111",
    "1111000011000110",
    "1111100010010100",
    "1111110110111100",
    "1111001111100100",
    "1110101110101001",
    "1110011001101111",
    "1110010011000001",
    "1110011000100010",
    "1110100101000000",
    "1110110010110110",
    "1110111110000100",
    "1111000101111011",
    "1111001110010111",
    "1111011100111111",
    "1111110101010100",
    "1111101001001001",
    "1111000011110001",
    "1110100010010010",
    "1110001011110101",
    "1110000100110001",
    "1110001100001010",
    "1110011100001111",
    "1110101110000010",
    "1110111100001010",
    "1111000100011101",
    "1111001000000100",
    "1111001001010001",
    "1111001100000010",
    "1111010101101100",
    "1111101001010100",
    "1111111001101101",
    "1111010111110001",
    "1110111000000001",
    "1110100001011001",
    "1110011000010001",
    "1110011101100001",
    "1110101101011001",
    "1111000001011001",
    "1111010011000101",
    "1111011111010110",
    "1111101000011101",
    "1111110011001101",
    "1111111100111010",
    "1111100111011000",
    "1111001111011110",
    "1110111011001001",
    "1110110000010010",
    "1110110001111110",
    "1110111110011110",
    "1111010000000010",
    "1111100000000111",
    "1111101010000001",
    "1111101101001110",
    "1111101101100101",
    "1111110000100011",
    "1111111010010010",
    "1111110100000011",
    "1111011101101101",
    "1111001000011011",
    "1110111010100000",
    "1110111000011011",
    "1111000010011101",
    "1111010100101111",
    "1111101001110010",
    "1111111100110100",
    "1111110101001000",
    "1111101101000110",
    "1111101010110111",
    "1111101101100001",
    "1111110011111001",
    "1111111101010010",
    "1111110110110101",
    "1111101001010010",
    "1111011010110010",
    "1111001100100110",
    "1111000000001101",
    "1110110110111110",
    "1110110001111011",
    "1110110001101100",
    "1110110110101000",
    "1111000000110101",
    "1111001111100100",
    "1111100001011110",
    "1111110100100100",
    "1111111001011110",
    "1111101010101101",
    "1111011111111000",
    "1111011000011101",
    "1111010010111001",
    "1111001101111010",
    "1111001001001001",
    "1111000101010011",
    "1111000011110001",
    "1111000101100111",
    "1111001011000111",
    "1111010011011101",
    "1111011100111000",
    "1111100101000000",
    "1111101001111100",
    "1111101010101110",
    "1111100111011000",
    "1111100000110011",
    "1111011000001100",
    "1111001110110000",
    "1111000101100101",
    "1110111101101011",
    "1110110111111001",
    "1110110101001110",
    "1110110110100010",
    "1110111100001111",
    "1111000101110110",
    "1111010010001010",
    "1111100000111011",
    "1111110011011010",
    "1111110101001100",
    "1111011001010000",
    "1110111011001010",
    "1110011111010010",
    "1110001010001100",
    "1101111111100110",
    "1110000000111000",
    "1110001011111000",
    "1110011100000111",
    "1110101100101011",
    "1110111011011101",
    "1111001010011011",
    "1111011100111010",
    "1111110100100110",
    "1111101111100011",
    "1111010011110001",
    "1110111101110000",
    "1110110010100001",
    "1110110100101111",
    "1111000100101001",
    "1111100000011010",
    "1111111011100001",
    "1111010100000110",
    "1110101110011100",
    "1110001111101001",
    "1101111100001110",
    "1101110110110100",
    "1101111111000111",
    "1110010001010111",
    "1110101001010101",
    "1111000101001000",
    "1111100100101001",
    "1111111000010000",
    "1111010011100001",
    "1110110000111001",
    "1110010100101110",
    "1110000011001000",
    "1101111111010001",
    "1110001000101000",
    "1110011011000001",
    "1110110000100110",
    "1111000011111001",
    "1111010010000101",
    "1111011100011100",
    "1111100111000001",
    "1111110110001001",
    "1111110100000000",
    "1111011001010110",
    "1110111110011011",
    "1110101000100111",
    "1110011100010110",
    "1110011011000010",
    "1110100010100110",
    "1110101111001000",
    "1110111100101010",
    "1111001000001000",
    "1111010000000101",
    "1111010100001010",
    "1111010100111100",
    "1111010100011000",
    "1111010101011010",
    "1111011011000010",
    "1111100110101111",
    "1111110111100111",
    "1111110101010011",
    "1111100100010101",
    "1111011001101111",
    "1111011000100101",
    "1111100001001000",
    "1111110000101011",
    "1111111100101001",
    "1111101010011001",
    "1111011010100110",
    "1111001101100110",
    "1111000011001010",
    "1110111011010100",
    "1110110110110111",
    "1110110111010000",
    "1110111101101011",
    "1111001001111001",
    "1111011010001011",
    "1111101011100101",
    "1111111011010001",
    "1111111000100110",
    "1111110000010100",
    "1111101010110010",
    "1111100110101111",
    "1111100011101100",
    "1111100010000101",
    "1111100011010010",
    "1111101000111000",
    "1111110011100010",
    "1111111101101100",
    "1111101101010010",
    "1111011110001100",
    "1111010011000011",
    "1111001101011110",
    "1111001101110011",
    "1111010011100001",
    "1111011101101000",
    "1111101011001010",
    "1111111011011000",
    "1111110010101011",
    "1111100000010111",
    "1111001111011100",
    "1111000010001011",
    "1110111010101010",
    "1110111010000110",
    "1111000000100001",
    "1111001100101101",
    "1111011100101011",
    "1111101110100000",
    "1111111111011101",
    "1111101110011110",
    "1111011111011001",
    "1111010010111101",
    "1111001001110101",
    "1111000100100000",
    "1111000011001011",
    "1111000101010011",
    "1111001010111000",
    "1111010101000011",
    "1111100101100100",
    "1111111101001011",
    "1111100101011101",
    "1111000110000000",
    "1110101001001110",
    "1110010011111110",
    "1110001001100101",
    "1110001010101101",
    "1110010110000001",
    "1110101001101111",
    "1111000100001101",
    "1111100011101001",
    "1111111010100101",
    "1111011010100000",
    "1111000000010001",
    "1110101111101110",
    "1110101011010100",
    "1110110010110001",
    "1111000011000000",
    "1111010111011011",
    "1111101011010101",
    "1111111011010010",
    "1111111001000110",
    "1111101110111100",
    "1111100010010000",
    "1111010000111011",
    "1110111100010100",
    "1110101000111100",
    "1110011100100110",
    "1110011100110101",
    "1110101100111111",
    "1111001100010110",
    "1111110110000001",
    "1111011101001010",
    "1110110100111001",
    "1110010111001001",
    "1110000111010011",
    "1110000101111110",
    "1110010000101100",
    "1110100011101110",
    "1110111100110010",
    "1111011011110101",
    "1111111110110110",
    "1111010100010111",
    "1110101000001100",
    "1101111111110101",
    "1101100000110000",
    "1101001111001100",
    "1101001100010011",
    "1101010101101010",
    "1101100110100111",
    "1101111001101101",
    "1110001010011000",
    "1110010110000110",
    "1110011100011110",
    "1110011110101011",
    "1110011110101001",
    "1110011110000101",
    "1110011101110010",
    "1110011110001101",
    "1110011111010001",
    "1110100001011010",
    "1110100111011011",
    "1110110100101001",
    "1111001010011000",
    "1111100110101100",
    "1111111011011011",
    "1111100001111001",
    "1111010001010111",
    "1111001100000101",
    "1111010000100011",
    "1111011001110000",
    "1111100001110110",
    "1111100100010111",
    "1111011111111011",
    "1111010110001011",
    "1111001010001111",
    "1110111111011110",
    "1110111001001011",
    "1110111010101010",
    "1111000110111111",
    "1111011111000100",
    "1111111111011110",
    "1111011001111010",
    "1110110110111111",
    "1110011101000111",
    "1110010000110011",
    "1110010010101110",
    "1110011111000010",
    "1110101111011111",
    "1110111110000010",
    "1111000111001000",
    "1111001010100010",
    "1111001001111100",
    "1111000111111111",
    "1111000110111100",
    "1111000111110001",
    "1111001010001100",
    "1111001101010110",
    "1111010000100100",
    "1111010011111110",
    "1111011000011101",
    "1111011110101001",
    "1111100110111011",
    "1111110001100100",
    "1111111110111000",
    "1111110001100111",
    "1111100001110001",
    "1111010100100010",
    "1111001100111101",
    "1111001101000101",
    "1111010101100101",
    "1111100101000011",
    "1111111000011000",
    "1111110100010000",
    "1111100100010111",
    "1111011010000111",
    "1111010110001000",
    "1111010111100111",
    "1111011100111100",
    "1111100100010010",
    "1111101100011000",
    "1111110100101011",
    "1111111101011100",
    "1111111000010111",
    "1111101100000011",
    "1111011101101001",
    "1111001101111111",
    "1110111110011001",
    "1110110000001100",
    "1110100100101001",
    "1110011100111000",
    "1110011001100010",
    "1110011010001110",
    "1110011101111011",
    "1110100010111110",
    "1110100111100101",
    "1110101010011001",
    "1110101010011110",
    "1110100111100010",
    "1110100010000101",
    "1110011010111111",
    "1110010011000101",
    "1110001010111100",
    "1110000010111001",
    "1101111011011000",
    "1101110101001011",
    "1101110001011110",
    "1101110001101011",
    "1101110110111110",
    "1110000001111011",
    "1110010010001010",
    "1110100110111110",
    "1110111111100110",
    "1111011011100000",
    "1111111001101110",
    "1111100111001101",
    "1111001001100111",
    "1110110000000111",
    "1110011101010001",
    "1110010010100010",
    "1110010000000000",
    "1110010100001010",
    "1110011100101000",
    "1110100110111011",
    "1110110001001111",
    "1110111100000001",
    "1111001010011000",
    "1111011111100110",
    "1111111100110100",
    "1111100000001010",
    "1110111100100110",
    "1110011110101001",
    "1110001011100101",
    "1110000101110100",
    "1110001011110101",
    "1110011001010011",
    "1110101001011000",
    "1110111000010000",
    "1111000100000101",
    "1111001100100110",
    "1111010010001010",
    "1111010101101001",
    "1111010111111100",
    "1111011001111010",
    "1111011100111000",
    "1111100010011010",
    "1111101011111110",
    "1111111010011100",
    "1111110010100011",
    "1111011101001010",
    "1111001000011010",
    "1110110111001011",
    "1110101010111010",
    "1110100011011000",
    "1110011111011100",
    "1110011101101101",
    "1110011100111111",
    "1110011101011011",
    "1110100000100111",
    "1110101000011011",
    "1110110101010010",
    "1111000100111100",
    "1111010010111101",
    "1111011010010001",
    "1111010111100000",
    "1111001010101010",
    "1110110111110010",
    "1110100101100010",
    "1110011010001100",
    "1110011001011000",
    "1110100010100110",
    "1110110010001011",
    "1111000011010111",
    "1111010001111110",
    "1111011100011110",
    "1111100101110111",
    "1111110011100101",
    "1111110110100111",
    "1111011000101010",
    "1110110110111111",
    "1110011000110100",
    "1110000100110110",
    "1101111111011110",
    "1110001000000100",
    "1110011001011110",
    "1110101101010110",
    "1110111110010111",
    "1111001010011110",
    "1111010100001110",
    "1111100000000111",
    "1111110001101111",
    "1111110110000100",
    "1111011011000110",
    "1111000011111001",
    "1110110110111100",
    "1110111001000001",
    "1111001010110010",
    "1111101000010011",
    "1111110100110110",
    "1111010011001101",
    "1110110111011000",
    "1110100011110011",
    "1110011001101000",
    "1110011000110101",
    "1110100000011001",
    "1110101110111000",
    "1111000010011101",
    "1111011000101100",
    "1111101110111010",
    "1111111101011010",
    "1111101110100001",
    "1111100101010011",
    "1111100001010000",
    "1111100001001000",
    "1111100011101100",
    "1111101000101101",
    "1111110000101000",
    "1111111011111010",
    "1111110101110001",
    "1111100101111110",
    "1111010111001001",
    "1111001011111111",
    "1111000110011101",
    "1111000111100010",
    "1111001111000111",
    "1111011100101010",
    "1111101111100000",
    "1111111001010101",
    "1111011111100001",
    "1111000101011101",
    "1110101101111111",
    "1110011100000010",
    "1110010010001010",
    "1110010001110110",
    "1110011010110000",
    "1110101010110101",
    "1110111110110101",
    "1111010011111001",
    "1111101000101111",
    "1111111101100111",
    "1111101100011001",
    "1111010100110100",
    "1110111100100001",
    "1110100110010000",
    "1110010101100111",
    "1110001101100011",
    "1110001111000000",
    "1110011000010101",
    "1110100101111001",
    "1110110011100110",
    "1110111110001111",
    "1111000100100111",
    "1111000111001011",
    "1111000111011111",
    "1111000111001011",
    "1111000111011010",
    "1111001000001100",
    "1111001000110101",
    "1111001000011101",
    "1111000110101101",
    "1111000100001000",
    "1111000001110001",
    "1111000000110110",
    "1111000010001000",
    "1111000101101111",
    "1111001011001111",
    "1111010001110001",
    "1111011001010101",
    "1111100100010010",
    "1111110101110000",
    "1111110001000000",
    "1111010001110011",
    "1110110001011110",
    "1110010110010010",
    "1110000101110111",
    "1110000011101010",
    "1110001110101110",
    "1110100010001011",
    "1110110111111110",
    "1111001010100110",
    "1111010111000001",
    "1111011100111000",
    "1111011101010100",
    "1111011011101010",
    "1111011101000010",
    "1111100101101110",
    "1111110111001101",
    "1111110000010011",
    "1111010101111100",
    "1110111111011001",
    "1110110001011001",
    "1110101110010110",
    "1110110101010111",
    "1111000010100100",
    "1111010001000111",
    "1111011100101010",
    "1111100011011111",
    "1111101000011000",
    "1111110000111011",
    "1111111110000111",
    "1111100011100010",
    "1111000011000000",
    "1110100011100100",
    "1110001100101010",
    "1110000011101111",
    "1110001001101011",
    "1110011001111010",
    "1110101101011100",
    "1110111110101011",
    "1111001100010001",
    "1111011001000110",
    "1111101000101101",
    "1111111101001111",
    "1111101010001010",
    "1111010010000000",
    "1111000000011111",
    "1110111011000111",
    "1111000100010000",
    "1111011010000111",
    "1111110111110001",
    "1111101000100010",
    "1111001011011110",
    "1110110011100010",
    "1110100010000011",
    "1110010111101111",
    "1110010100110011",
    "1110011001101010",
    "1110100111011010",
    "1110111110100001",
    "1111011101101000",
    "1111111111001011",
    "1111011101101110",
    "1111000011100010",
    "1110110100100010",
    "1110110001111110",
    "1110111010100011",
    "1111001011001001",
    "1111100000100011",
    "1111111000100001",
    "1111101110000001",
    "1111010011111001",
    "1110111010100110",
    "1110100100011101",
    "1110010100000110",
    "1110001011100011",
    "1110001011110000",
    "1110010100011010",
    "1110100100101001",
    "1110111011010011",
    "1111010110110010",
    "1111110101011101",
    "1111101010011100",
    "1111001011001110",
    "1110101111100100",
    "1110011010001110",
    "1110001101000000",
    "1110001000001000",
    "1110001001111101",
    "1110010000001111",
    "1110011001000100",
    "1110100011110110",
    "1110110001001111",
    "1111000010001011",
    "1111010110111100",
    "1111101110000111",
    "1111111011000110",
    "1111101000001000",
    "1111011011101111",
    "1111010110110010",
    "1111011000000100",
    "1111011100111100",
    "1111100010100001",
    "1111100110110111",
    "1111101001011000",
    "1111101010100110",
    "1111101011100101",
    "1111101101001011",
    "1111101111010001",
    "1111110000101011",
    "1111101111100001",
    "1111101010001110",
    "1111100000001000",
    "1111010001101100",
    "1111000000011111",
    "1110101110111000",
    "1110011111101001",
    "1110010101011010",
    "1110010001111001",
    "1110010101101010",
    "1110100001000111",
    "1110110101011011",
    "1111010011001101",
    "1111111000110011",
    "1111011101111111",
    "1110110111011111",
    "1110011001110101",
    "1110001001100011",
    "1110001000001011",
    "1110010010111110",
    "1110100100001110",
    "1110110101111100",
    "1111000011101100",
    "1111001011110010",
    "1111001111000100",
    "1111001111011001",
    "1111001111011001",
    "1111010011011111",
    "1111100000001000",
    "1111110111001000",
    "1111101000111111",
    "1111000101011000",
    "1110100100101110",
    "1110001100110000",
    "1110000001011010",
    "1110000011000001",
    "1110001101110010",
    "1110011011111101",
    "1110101000001110",
    "1110101111001111",
    "1110110001000011",
    "1110101111010001",
    "1110101100110101",
    "1110101111000000",
    "1110111010011011",
    "1111010000101110",
    "1111110000000011",
    "1111101101000001",
    "1111001101010010",
    "1110110110001011",
    "1110101011001111",
    "1110101101000000",
    "1110111001000010",
    "1111001011110101",
    "1111100001100001",
    "1111110111000011",
    "1111110101010100",
    "1111100101011111",
    "1111011011000110",
    "1111010111001001",
    "1111011010001111",
    "1111100011101001",
    "1111110001010110",
    "1111111110111110",
    "1111101111110111",
    "1111100011100100",
    "1111011011110000",
    "1111011001010110",
    "1111011100011110",
    "1111100100111100",
    "1111110010101110",
    "1111111010110101",
    "1111100101101111",
    "1111010000100110",
    "1110111110001010",
    "1110110000011111",
    "1110101000100111",
    "1110100110101010",
    "1110101001111100",
    "1110110001000011",
    "1110111010011110",
    "1111000101101001",
    "1111010011011100",
    "1111100101011000",
    "1111111100011110",
    "1111100111111100",
    "1111001010100000",
    "1110101111010010",
    "1110011010111010",
    "1110010001001000",
    "1110010011011010",
    "1110100000101011",
    "1110110101101100",
    "1111001110010100",
    "1111100110001110",
    "1111111001100000",
    "1111111010111100",
    "1111111001000101",
    "1111111111000011",
    "1111101111110000",
    "1111011100110011",
    "1111001010101000",
    "1110111100111101",
    "1110110101111001",
    "1110110101010011",
    "1110111000111110",
    "1110111101101110",
    "1111000001000111",
    "1111000010001010",
    "1111000001101100",
    "1111000010101100",
    "1111001001110101",
    "1111011010100101",
    "1111110101011010",
    "1111101001000101",
    "1111000111010000",
    "1110101011100110",
    "1110011011001111",
    "1110011000001110",
    "1110100000011010",
    "1110101111001111",
    "1111000000000000",
    "1111001111001101",
    "1111011011110111",
    "1111100110010110",
    "1111110000000110",
    "1111111100000011",
    "1111110010111110",
    "1111011100100101",
    "1111000010110100",
    "1110101010001111",
    "1110010111111100",
    "1110001111011110",
    "1110010010010000",
    "1110011110101011",
    "1110110001010100",
    "1111000111001110",
    "1111011111000000",
    "1111111000011001",
    "1111101100100111",
    "1111010001010100",
    "1110111000100000",
    "1110100101100101",
    "1110011100001001",
    "1110011110000000",
    "1110101001111101",
    "1110111100111010",
    "1111010100101001",
    "1111110000001111",
    "1111110000111111",
    "1111010000010111",
    "1110110000101100",
    "1110010110000011",
    "1110000100110111",
    "1110000000011001",
    "1110001000001100",
    "1110010111111100",
    "1110101001101010",
    "1110111000000001",
    "1111000000010101",
    "1111000011000110",
    "1111000011011010",
    "1111000110001001",
    "1111001111111000",
    "1111100010000110",
    "1111111010111111",
    "1111101001111101",
    "1111010010010100",
    "1111000010010010",
    "1110111011100011",
    "1110111100111000",
    "1111000011001000",
    "1111001011000001",
    "1111010010010000",
    "1111011000001001",
    "1111011101100000",
    "1111100011111000",
    "1111101100100000",
    "1111110111011010",
    "1111111100101010",
    "1111110010001011",
    "1111101011011110",
    "1111101010010111",
    "1111101111011010",
    "1111111001111011",
    "1111110111100010",
    "1111100110101000",
    "1111010101000101",
    "1111000100110110",
    "1110110111111001",
    "1110101111101100",
    "1110101100101110",
    "1110101110011011",
    "1110110011101111",
    "1110111011100001",
    "1111000100101100",
    "1111001110101011",
    "1111011001001001",
    "1111100100001011",
    "1111101111111110",
    "1111111100111101",
    "1111110100101011",
    "1111100101100101",
    "1111010111001101",
    "1111001011010110",
    "1111000011010101",
    "1110111111100100",
    "1110111111100011",
    "1111000010001011",
    "1111000110001011",
    "1111001010101010",
    "1111001111010111",
    "1111010100011100",
    "1111011010000110",
    "1111100000000010",
    "1111100101101111",
    "1111101010010010",
    "1111101100110001",
    "1111101100101010",
    "1111101010010101",
    "1111100110111100",
    "1111100100000011",
    "1111100011000000",
    "1111100100101110",
    "1111101001100000",
    "1111110001001101",
    "1111111011010011",
    "1111111000111111",
    "1111101100110001",
    "1111100001000000",
    "1111010110100000",
    "1111001101110101",
    "1111000110111001",
    "1111000001010101",
    "1110111100101011",
    "1110111000011101",
    "1110110100100010",
    "1110110001001010",
    "1110101110101110",
    "1110101101111000",
    "1110101111001101",
    "1110110011011000",
    "1110111011011000",
    "1111001000000100",
    "1111011001010011",
    "1111101101100011",
    "1111111101111001",
    "1111101100100010",
    "1111100001010111",
    "1111011110001100",
    "1111100010101111",
    "1111101100110000",
    "1111111000111110",
    "1111111011110000",
    "1111110011110110",
    "1111110000011000",
    "1111110001011110",
    "1111110110101001",
    "1111111111001111",
    "1111110101010010",
    "1111100111100110",
    "1111011000011000",
    "1111001000100111",
    "1110111001010101",
    "1110101011110011",
    "1110100001010100",
    "1110011010110101",
    "1110011000110010",
    "1110011010111000",
    "1110100000010101",
    "1110100111111001",
    "1110110000000111",
    "1110110111100111",
    "1110111110001100",
    "1111000101111110",
    "1111010010000110",
    "1111100100100101",
    "1111111100101010",
    "1111101001100111",
    "1111010100011101",
    "1111001010000010",
    "1111001110110011",
    "1111100011001101",
    "1111111100110100",
    "1111011000010000",
    "1110110110110110",
    "1110011110110101",
    "1110010011011101",
    "1110010101010011",
    "1110100010100110",
    "1110111000010110",
    "1111010011100010",
    "1111110001011011",
    "1111110000011001",
    "1111010100001000",
    "1110111011111010",
    "1110101001101101",
    "1110011110110001",
    "1110011011000110",
    "1110011101010010",
    "1110100011011111",
    "1110101011100011",
    "1110110011101111",
    "1110111010110100",
    "1111000000010111",
    "1111000101001011",
    "1111001011001110",
    "1111010101001110",
    "1111100101011101",
    "1111111100011110",
    "1111100111100101",
    "1111001010110111",
    "1110110010011100",
    "1110100010111000",
    "1110011110101101",
    "1110100101100010",
    "1110110100010000",
    "1111000110010011",
    "1111010110111111",
    "1111100010110011",
    "1111101000000111",
    "1111100111000101",
    "1111100001001100",
    "1111011000010110",
    "1111001110011110",
    "1111000101011000",
    "1110111111010110",
    "1110111110101101",
    "1111000101010011",
    "1111010011010010",
    "1111100110100111",
    "1111111011011011",
    "1111110010101011",
    "1111100111011011",
    "1111100100100010",
    "1111101001010010",
    "1111110010110110",
    "1111111101100000",
    "1111111010001101",
    "1111110110101010",
    "1111111000111011",
    "1111111111000010",
    "1111110010010010",
    "1111100010001101",
    "1111010000010101",
    "1110111110011100",
    "1110101110011111",
    "1110100010100111",
    "1110011100100110",
    "1110011101101101",
    "1110100111000001",
    "1110111001011000",
    "1111010100010010",
    "1111110101001001",
    "1111101000011011",
    "1111001001111100",
    "1110110100001110",
    "1110101010001110",
    "1110101011110000",
    "1110110101010101",
    "1111000001101100",
    "1111001100010100",
    "1111010011101010",
    "1111011001101101",
    "1111100010000110",
    "1111110000000111",
    "1111111011000011",
    "1111100001001101",
    "1111000110001101",
    "1110101110110101",
    "1110011110111011",
    "1110011000010011",
    "1110011010111101",
    "1110100110001101",
    "1110111001010001",
    "1111010011010011",
    "1111110010001010",
    "1111101101111010",
    "1111010001101011",
    "1110111101011110",
    "1110110100001000",
    "1110110101111001",
    "1111000000101100",
    "1111010001010010",
    "1111100100111011",
    "1111111010100010",
    "1111101101110001",
    "1111010100001101",
    "1110111010010001",
    "1110100011000000",
    "1110010010001000",
    "1110001010100101",
    "1110001101010001",
    "1110011000100010",
    "1110101001010011",
    "1110111101100001",
    "1111010100111001",
    "1111110000000100",
    "1111110001001111",
    "1111010001100010",
    "1110110101010101",
    "1110100001110110",
    "1110011011001001",
    "1110100001111110",
    "1110110011010010",
    "1111001001100011",
    "1111011111000100",
    "1111101111111010",
    "1111111011011101",
    "1111111011000101",
    "1111101110110001",
    "1111011100001111",
    "1111000100010101",
    "1110101100010011",
    "1110011011110101",
    "1110011001101101",
    "1110101001001001",
    "1111000111111110",
    "1111101111000010",
    "1111101010100000",
    "1111001100010001",
    "1110111010100000",
    "1110110101101100",
    "1110111100001010",
    "1111001011110010",
    "1111100010100100",
    "1111111110110111",
    "1111100001010111",
    "1111000001011010",
    "1110100101010000",
    "1110010001000010",
    "1110000111101101",
    "1110001001101111",
    "1110010100100010",
    "1110100011100010",
    "1110110010000101",
    "1110111101000100",
    "1111000011010111",
    "1111000101011011",
    "1111000100100010",
    "1111000010001000",
    "1110111111010001",
    "1110111100100011",
    "1110111010011101",
    "1110111010011101",
    "1110111111101110",
    "1111001100111101",
    "1111100010010100",
    "1111111100100111",
    "1111101010000000",
    "1111011000000001",
    "1111010010001111",
    "1111011010100000",
    "1111101110011111",
    "1111110111001000",
    "1111011100010111",
    "1111000110000011",
    "1110110110110001",
    "1110101111000000",
    "1110101110010001",
    "1110110011000110",
    "1110111100000101",
    "1111001000100000",
    "1111011000010011",
    "1111101011110000",
    "1111111101010111",
    "1111100100100111",
    "1111001100100011",
    "1110110111111001",
    "1110101000011110",
    "1110011110111011",
    "1110011010111100",
    "1110011011001110",
    "1110011110000100",
    "1110100001110001",
    "1110100101011010",
    "1110101000110100",
    "1110101100101000",
    "1110110011011100",
    "1111000001001010",
    "1111011000001100",
    "1111110111100101",
    "1111100101001101",
    "1111000101011000",
    "1110101111111000",
    "1110101001111100",
    "1110110101011101",
    "1111001111111000",
    "1111110011010011",
    "1111100111101111",
    "1111001000110010",
    "1110110100111001",
    "1110101110100100",
    "1110110110000100",
    "1111001001101010",
    "1111100110010011",
    "1111110111101011",
    "1111010100110011",
    "1110110101001101",
    "1110011100011110",
    "1110001100111111",
    "1110000111100101",
    "1110001011000111",
    "1110010100111011",
    "1110100010011111",
    "1110110011001010",
    "1111001000000110",
    "1111100010100100",
    "1111111101011011",
    "1111011010001110",
    "1110110111011111",
    "1110011001010001",
    "1110000010111110",
    "1101110110011101",
    "1101110011110110",
    "1101111010011001",
    "1110001001100111",
    "1110100001010010",
    "1111000000111011",
    "1111100110100010",
    "1111110001101100",
    "1111001100111101",
    "1110110000101011",
    "1110100000110011",
    "1110011110011110",
    "1110100111110100",
    "1110111000110111",
    "1111001100111101",
    "1111100000010101",
    "1111110000111010",
    "1111111110011100",
    "1111110110001001",
    "1111101100100000",
    "1111100101100101",
    "1111100011011111",
    "1111101000100101",
    "1111110110010000",
    "1111110100011001",
    "1111011010111111",
    "1111000010110011",
    "1110110000110110",
    "1110101000000100",
    "1110101000100111",
    "1110110000000010",
    "1110111010110101",
    "1111000101101100",
    "1111001110111011",
    "1111011001010000",
    "1111101010000010",
    "1111111011000010",
    "1111010110011010",
    "1110101101001010",
    "1110000111011111",
    "1101101100111111",
    "1101100010101110",
    "1101101000111001",
    "1101111010010110",
    "1110001111111111",
    "1110100011101001",
    "1110110001111000",
    "1110111010101010",
    "1111000000111110",
    "1111001010010110",
    "1111011011110010",
    "1111110110001011",
    "1111101010000110",
    "1111001011111010",
    "1110110110010101",
    "1110101110000111",
    "1110110100000011",
    "1111000100001010",
    "1111010111111100",
    "1111101001101000",
    "1111110101011010",
    "1111111010001101",
    "1111111001011100",
    "1111110101110100",
    "1111110011110001",
    "1111111000011011",
    "1111111001000010",
    "1111100000110011",
    "1111000010011101",
    "1110100100001110",
    "1110001100010001",
    "1101111110111000",
    "1101111101100110",
    "1110000110110111",
    "1110010111011000",
    "1110101011001110",
    "1110111111000111",
    "1111010001011010",
    "1111100001111101",
    "1111110000110111",
    "1111111110000100",
    "1111110111010110",
    "1111110001000010",
    "1111110000001100",
    "1111110101010000",
    "1111111111111000",
    "1111110000001111",
    "1111011101011110",
    "1111001001101000",
    "1110110110110010",
    "1110100110111011",
    "1110011011110010",
    "1110010110100000",
    "1110010111000100",
    "1110011100010100",
    "1110100100011111",
    "1110101110000000",
    "1110111000100010",
    "1111000101001101",
    "1111010101100000",
    "1111101001110000",
    "1111111111110000",
    "1111101010101101",
    "1111011011100000",
    "1111010110010101",
    "1111011110010100",
    "1111110011101101",
    "1111101100010001",
    "1111000110100010",
    "1110100000110000",
    "1110000000100001",
    "1101101010010100",
    "1101100000110110",
    "1101100100011101",
    "1101110011001000",
    "1110001001101000",
    "1110100100010010",
    "1111000000000111",
    "1111011011001111",
    "1111110100111001",
    "1111110011001010",
    "1111011101001010",
    "1111001001110100",
    "1110111010101000",
    "1110110001100111",
    "1110110000010111",
    "1110110111000110",
    "1111000100100000",
    "1111010101110100",
    "1111100111100110",
    "1111110110111110",
    "1111111101110000",
    "1111110110111111",
    "1111110100000011",
    "1111110011110100",
    "1111110101100011",
    "1111111000111000",
    "1111111101101110",
    "1111111100011100",
    "1111110110110101",
    "1111110011001011",
    "1111110011001111",
    "1111111000010011",
    "1111111101001111",
    "1111101110001100",
    "1111011100010001",
    "1111001001100111",
    "1110111000010001",
    "1110101001111010",
    "1110011111101011",
    "1110011010001111",
    "1110011001111010",
    "1110011110100001",
    "1110100111011111",
    "1110110011101100",
    "1111000001111000",
    "1111010000100111",
    "1111011111100011",
    "1111110000000010",
    "1111111011010011",
    "1111100000110011",
    "1111000000101011",
    "1110011110000010",
    "1101111101111111",
    "1101100101111100",
    "1101011001111111",
    "1101011010110101",
    "1101100101110001",
    "1101110101111110",
    "1110000110011010",
    "1110010011011101",
    "1110011100010011",
    "1110100011010101",
    "1110101100110011",
    "1110111100000001",
    "1111010001000011",
    "1111101000100011",
    "1111111101000101",
    "1111110110100111",
    "1111110101111001",
    "1111111111011110",
    "1111101101000011",
    "1111010111100011",
    "1111000011010111",
    "1110110011011000",
    "1110101000111001",
    "1110100011111000",
    "1110100011011000",
    "1110100101110010",
    "1110101001011011",
    "1110101100011011",
    "1110101101001001",
    "1110101010011110",
    "1110100100001010",
    "1110011011000110",
    "1110010001001111",
    "1110001001000110",
    "1110000101011010",
    "1110001001001001",
    "1110010110000011",
    "1110101011100001",
    "1111000110101010",
    "1111100010110011",
    "1111111011001000",
    "1111110100000010",
    "1111101100100001",
    "1111101101011000",
    "1111110011010001",
    "1111111010000011",
    "1111111110010001",
    "1111111110010011",
    "1111111010011001",
    "1111110100011001",
    "1111101111011010",
    "1111101110011111",
    "1111110011000010",
    "1111111100001011",
    "1111111000111111",
    "1111110000100100",
    "1111101110001000",
    "1111110011101101",
    "1111111110110101",
    "1111101011111000",
    "1111010110111011",
    "1111000011111001",
    "1110110110001000",
    "1110101111100001",
    "1110110000101001",
    "1110111001000010",
    "1111000111111110",
    "1111011100110011",
    "1111110111001000",
    "1111101001110100",
    "1111000111110111",
    "1110100110001011",
    "1110001001001100",
    "1101110101011000",
    "1101101101100110",
    "1101110010000101",
    "1110000000011010",
    "1110010100100010",
    "1110101010000110",
    "1110111110011100",
    "1111010001100111",
    "1111100101010010",
    "1111111010110110",
    "1111101101110001",
    "1111010111001110",
    "1111000101011101",
    "1110111100001001",
    "1110111100110000",
    "1111000101011000",
    "1111010001101100",
    "1111011100110011",
    "1111100011000000",
    "1111100011000011",
    "1111011110000100",
    "1111010110101000",
    "1111001111110011",
    "1111001011101011",
    "1111001010100110",
    "1111001011100000",
    "1111001100100001",
    "1111001011111010",
    "1111001000111010",
    "1111000011111100",
    "1110111110011110",
    "1110111010010110",
    "1110111001010011",
    "1110111101111000",
    "1111001011110010",
    "1111100101001101",
    "1111110110111001",
    "1111001101011011",
    "1110100101110001",
    "1110000111010110",
    "1101110111011010",
    "1101110111100000",
    "1110000100010101",
    "1110010111101010",
    "1110101011001110",
    "1110111010100010",
    "1111000100001010",
    "1111001001001001",
    "1111001011011011",
    "1111001101001110",
    "1111001111100110",
    "1111010010111000",
    "1111011000111001",
    "1111100100000101",
    "1111110101101111",
    "1111110010110011",
    "1111011001010000",
    "1111000011001101",
    "1110110110100100",
    "1110110111101010",
    "1111000110101000",
    "1111011111010010",
    "1111111011011101",
    "1111101011000110",
    "1111011000111100",
    "1111001111111111",
    "1111010000010001",
    "1111011000011000",
    "1111100110000100",
    "1111110111100000",
    "1111110101000110",
    "1111100001101110",
    "1111010000011010",
    "1111000011100001",
    "1110111101000000",
    "1110111101111010",
    "1111000101101010",
    "1111010010001010",
    "1111100000100011",
    "1111101110011011",
    "1111111010010011",
    "1111111100010111",
    "1111110101010100",
    "1111101111110011",
    "1111101010110111",
    "1111100101100101",
    "1111011111001100",
    "1111010111100000",
    "1111001110110110",
    "1111000110011101",
    "1111000000000010",
    "1110111101001100",
    "1110111110111011",
    "1111000101010101",
    "1111001111011111",
    "1111011101001111",
    "1111101111101011",
    "1111111000100000",
    "1111011100010100",
    "1110111110111000",
    "1110100101010111",
    "1110010101000011",
    "1110010001111001",
    "1110011100101000",
    "1110110001010000",
    "1111001000111111",
    "1111011100110111",
    "1111100111111101",
    "1111101001010100",
    "1111100011010000",
    "1111011011100110",
    "1111011010011000",
    "1111100101001110",
    "1111111100101110",
    "1111100011110100",
    "1111000100101100",
    "1110101110000010",
    "1110100101011011",
    "1110101100000111",
    "1110111110010111",
    "1111010110100010",
    "1111110000000111",
    "1111110111000011",
    "1111011111001010",
    "1111000111111111",
    "1110110010110001",
    "1110100001101110",
    "1110010111101111",
    "1110010111011010",
    "1110100001000010",
    "1110110010001111",
    "1111000111000011",
    "1111011011000001",
    "1111101010101111",
    "1111110100101100",
    "1111111000111110",
    "1111111000001110",
    "1111110011000110",
    "1111101001111111",
    "1111011101111011",
    "1111010001000011",
    "1111000101111011",
    "1110111111010010",
    "1110111111011001",
    "1111000111011000",
    "1111010111000011",
    "1111101100100010",
    "1111111011001010",
    "1111100011011000",
    "1111001110110101",
    "1110111111010100",
    "1110110101011011",
    "1110110000100100",
    "1110101111010100",
    "1110101111111010",
    "1110110001001101",
    "1110110011010111",
    "1110110111111100",
    "1111000001010101",
    "1111010001011111",
    "1111101000110101",
    "1111111010010100",
    "1111011011101111",
    "1110111111111010",
    "1110101010111010",
    "1110011111000100",
    "1110011100000111",
    "1110100000001100",
    "1110101000011101",
    "1110110010001101",
    "1110111011011000",
    "1111000010110011",
    "1111001000110111",
    "1111001111011001",
    "1111011000101010",
    "1111100110001110",
    "1111110111111101",
    "1111110100000000",
    "1111100000101011",
    "1111010001000101",
    "1111000111100111",
    "1111000100110110",
    "1111000111100101",
    "1111001101100000",
    "1111010011111011",
    "1111011001101111",
    "1111100000010100",
    "1111101010010011",
    "1111111001101011",
    "1111110001111000",
    "1111011100000010",
    "1111001010011011",
    "1111000011000011",
    "1111001001111101",
    "1111011110110110",
    "1111111101001000",
    "1111100010001000",
    "1111000110001011",
    "1110110100001000",
    "1110101110011011",
    "1110110101010010",
    "1111000111010110",
    "1111100010001010",
    "1111111101001101",
    "1111011010001110",
    "1110111000100000",
    "1110011011101111",
    "1110000111001110",
    "1101111101001010",
    "1101111101100011",
    "1110000110001110",
    "1110010011110011",
    "1110100011111100",
    "1110110110110111",
    "1111001110001101",
    "1111101011001011",
    "1111110011000110",
    "1111010000001000",
    "1110110000110101",
    "1110011001111001",
    "1110001110010111",
    "1110001101110101",
    "1110010100111001",
    "1110011111001000",
    "1110101000111111",
    "1110110000111000",
    "1110110111000011",
    "1110111100100101",
    "1111000010110001",
    "1111001010100010",
    "1111010100100111",
    "1111100010100001",
    "1111110101011010",
    "1111110010111010",
    "1111011000111001",
    "1111000001001000",
    "1110110001011110",
    "1110101111001000",
    "1110111100110010",
    "1111011000010101",
    "1111111011100101",
    "1111100001001010",
    "1111000100110001",
    "1110110011000011",
    "1110101100100000",
    "1110101110111010",
    "1110110110110001",
    "1111000001001010",
    "1111001101111000",
    "1111011110100011",
    "1111110100111001",
    "1111101111001111",
    "1111010000111110",
    "1110110101001001",
    "1110100000101110",
    "1110010110111111",
    "1110011000010001",
    "1110100001111001",
    "1110101111100001",
    "1110111100111100",
    "1111000111100000",
    "1111001111010111",
    "1111010111011000",
    "1111100011010101",
    "1111110101101010",
    "1111110010011010",
    "1111011001000110",
    "1111000100001010",
    "1110111001001001",
    "1110111011110000",
    "1111001100100011",
    "1111101001010011",
    "1111110010000001",
    "1111001010011110",
    "1110100101001001",
    "1110000110110110",
    "1101110011010010",
    "1101101100001111",
    "1101110001000011",
    "1101111111011110",
    "1110010100110111",
    "1110101111011010",
    "1111001101101110",
    "1111101110010010",
    "1111110001001101",
    "1111010011101100",
    "1110111011110000",
    "1110101011011001",
    "1110100011100001",
    "1110100011011111",
    "1110101001001001",
    "1110110001010100",
    "1110111001000100",
    "1110111110101011",
    "1111000010100010",
    "1111000111001000",
    "1111001111110110",
    "1111011111010100",
    "1111110101101111",
    "1111101111100000",
    "1111010101001011",
    "1111000000010101",
    "1110110100101100",
    "1110110011100100",
    "1110111011100101",
    "1111001001010001",
    "1111011000010101",
    "1111100100110001",
    "1111101011111010",
    "1111101100110010",
    "1111100111101110",
    "1111011101111101",
    "1111010000111110",
    "1111000010010111",
    "1110110011101100",
    "1110100110011010",
    "1110011011110010",
    "1110010100110011",
    "1110010010000000",
    "1110010011011101",
    "1110011000110010",
    "1110100001000011",
    "1110101011000010",
    "1110110101010011",
    "1110111110100110",
    "1111000110001000",
    "1111001100000101",
    "1111010011000110",
    "1111011111011110",
    "1111110100100001",
    "1111101101011101",
    "1111001010001100",
    "1110101000000100",
    "1110001110010010",
    "1110000011001111",
    "1110001010100101",
    "1110100011010111",
    "1111001000011010",
    "1111110010000010",
    "1111100111100111",
    "1111001010011101",
    "1110111001100011",
    "1110110101001101",
    "1110111011000010",
    "1111000111111100",
    "1111011001110111",
    "1111101111110011",
    "1111110110101101",
    "1111011011000100",
    "1111000000010100",
    "1110101010011011",
    "1110011101000111",
    "1110011010011011",
    "1110100010001000",
    "1110110001110100",
    "1111000101110100",
    "1111011001111111",
    "1111101011001000",
    "1111110111101101",
    "1111111111111101",
    "1111111010100101",
    "1111110110001011",
    "1111110001010101",
    "1111101011011100",
    "1111100100100111",
    "1111011101110111",
    "1111011000101010",
    "1111010110011011",
    "1111011000001001",
    "1111011110000010",
    "1111100111111101",
    "1111110101101010",
    "1111111001001010",
    "1111100101010010",
    "1111010000000000",
    "1110111011011001",
    "1110101010000001",
    "1110011110010001",
    "1110011001100011",
    "1110011011100101",
    "1110100010001111",
    "1110101010101000",
    "1110110001111110",
    "1110110110011101",
    "1110110111011011",
    "1110110101000110",
    "1110110000101001",
    "1110101100001010",
    "1110101010011110",
    "1110101110000111",
    "1110111000001001",
    "1111000111011101",
    "1111011001000110",
    "1111101000111111",
    "1111110011000110",
    "1111110100111010",
    "1111101110011011",
    "1111100010001010",
    "1111010011111110",
    "1111000111101111",
    "1111000000001111",
    "1110111110111011",
    "1111000100000000",
    "1111001110111010",
    "1111011110100110",
    "1111110001110011",
    "1111111000111100",
    "1111100011110110",
    "1111010001011010",
    "1111000100001000",
    "1110111101100110",
    "1110111101111011",
    "1111000011110110",
    "1111001101001001",
    "1111010111011000",
    "1111100000101110",
    "1111101000011001",
    "1111101110111000",
    "1111110101011010",
    "1111111101001011",
    "1111111001010111",
    "1111101111000011",
    "1111100101001110",
    "1111011101010111",
    "1111011000010000",
    "1111010101100111",
    "1111010100100100",
    "1111010100001000",
    "1111010011110100",
    "1111010011100100",
    "1111010011101010",
    "1111010100010010",
    "1111010100111100",
    "1111010100011101",
    "1111010001100010",
    "1111001011011001",
    "1111000010011001",
    "1110110111110101",
    "1110101101100100",
    "1110100101010000",
    "1110011111111101",
    "1110011101110101",
    "1110011110010110",
    "1110100000101011",
    "1110100100000101",
    "1110101000001011",
    "1110101100101101",
    "1110110001011010",
    "1110110101111100",
    "1110111010000010",
    "1110111101100100",
    "1111000001001111",
    "1111000111010000",
    "1111010010010111",
    "1111100011111110",
    "1111111010111000",
    "1111101101000000",
    "1111011001110101",
    "1111010001100110",
    "1111011000011000",
    "1111101110010100",
    "1111110000111110",
    "1111001100101011",
    "1110101100100001",
    "1110010110101000",
    "1110001110011110",
    "1110010101111110",
    "1110101101001111",
    "1111010001110110",
    "1111111111000100",
    "1111010001110110",
    "1110101000011000",
    "1110001010101011",
    "1101111100010111",
    "1101111101001010",
    "1110001000110010",
    "1110011000101100",
    "1110100110100111",
    "1110101110110110",
    "1110110001000010",
    "1110101111010001",
    "1110101100100101",
    "1110101100010100",
    "1110110010011100",
    "1111000010000010",
    "1111011011110000",
    "1111111100110111",
    "1111100000000111",
    "1111000001101001",
    "1110101100111000",
    "1110100101000110",
    "1110101001111101",
    "1110110111011010",
    "1111000111101000",
    "1111010101010111",
    "1111011101100011",
    "1111011111111000",
    "1111011101011100",
    "1111011000010011",
    "1111010010100001",
    "1111001101010110",
    "1111001010001001",
    "1111001011010001",
    "1111010010111011",
    "1111100010010101",
    "1111111000110110",
    "1111101100100011",
    "1111010010110110",
    "1110111111011100",
    "1110110110011010",
    "1110111000101100",
    "1111000100011010",
    "1111010110000110",
    "1111101001100111",
    "1111111011001111",
    "1111110111101011",
    "1111110000110111",
    "1111110000100011",
    "1111110110000000",
    "1111111111111100",
    "1111110010110101",
    "1111100011101110",
    "1111010010111011",
    "1111000000110001",
    "1110101110010110",
    "1110011101110000",
    "1110010001011111",
    "1110001011001110",
    "1110001011100000",
    "1110010001011010",
    "1110011011010110",
    "1110101000000100",
    "1110110111010000",
    "1111001000111111",
    "1111011101001001",
    "1111110010110101",
    "1111110111111000",
    "1111100101011101",
    "1111011000001001",
    "1111010001001000",
    "1111010000010010",
    "1111010100010011",
    "1111011011101000",
    "1111100100111110",
    "1111101111100010",
    "1111111010100110",
    "1111111010010111",
    "1111101111111001",
    "1111100110011100",
    "1111011110100110",
    "1111011001000001",
    "1111010110000011",
    "1111010101110001",
    "1111010111100101",
    "1111011010101111",
    "1111011110001100",
    "1111100000111001",
    "1111100010000000",
    "1111100000111101",
    "1111011101101110",
    "1111011000111111",
    "1111010011101111",
    "1111001111000010",
    "1111001011101101",
    "1111001010001011",
    "1111001010100011",
    "1111001100111000",
    "1111010000110000",
    "1111010101100000",
    "1111011010010001",
    "1111011110001100",
    "1111100000110110",
    "1111100010011001",
    "1111100011011010",
    "1111100100101010",
    "1111100110100100",
    "1111101000110110",
    "1111101010110110",
    "1111101011110010",
    "1111101011001000",
    "1111101000110011",
    "1111100101010010",
    "1111100001000010",
    "1111011100001010",
    "1111010110001000",
    "1111001101111000",
    "1111000010101100",
    "1110110100100100",
    "1110100100100111",
    "1110010101000110",
    "1110001000110101",
    "1110000010101001",
    "1110000100100101",
    "1110010000000101",
    "1110100101010111",
    "1111000011000001",
    "1111100101101110",
    "1111110111010111",
    "1111011001011000",
    "1111000100101010",
    "1110111011110111",
    "1110111111110000",
    "1111001111011111",
    "1111101000110010",
    "1111110111110100",
    "1111010110110001",
    "1110111000100011",
    "1110100001010010",
    "1110010011101010",
    "1110010000100001",
    "1110010110100101",
    "1110100011000110",
    "1110110011000101",
    "1111000100101111",
    "1111010111011011",
    "1111101010111101",
    "1111111110110000",
    "1111101110010001",
    "1111011110000000",
    "1111010010011100",
    "1111001101000111",
    "1111001110000100",
    "1111010011011111",
    "1111011010011110",
    "1111100000000000",
    "1111100010000110",
    "1111100000011111",
    "1111011100010100",
    "1111010111011011",
    "1111010011101001",
    "1111010010100100",
    "1111010101110110",
    "1111011110111111",
    "1111101110010110",
    "1111111101100100",
    "1111101000010011",
    "1111010110010011",
    "1111001011101011",
    "1111001010110111",
    "1111010011100001",
    "1111100010011010",
    "1111110010110000",
    "1111111111111000",
    "1111111000011001",
    "1111110110100101",
    "1111110110100000",
    "1111110010101011",
    "1111100111001101",
    "1111010011110110",
    "1110111100100110",
    "1110100111111010",
    "1110011100000001",
    "1110011101100001",
    "1110101101101000",
    "1111001010001100",
    "1111101110110100",
    "1111101010000000",
    "1111000101101100",
    "1110101000100000",
    "1110010101011111",
    "1110001101100011",
    "1110001111011111",
    "1110011000100000",
    "1110100101000001",
    "1110110001111000",
    "1110111101001100",
    "1111000111100000",
    "1111010011110011",
    "1111100101000110",
    "1111111100110011",
    "1111100110110000",
    "1111001010011000",
    "1110110100010111",
    "1110101010011101",
    "1110101111101001",
    "1111000010010101",
    "1111011101001100",
    "1111111001011101",
    "1111101111000100",
    "1111100000011111",
    "1111011100101110",
    "1111100100000000",
    "1111110100110101",
    "1111110011010001",
    "1111010111100010",
    "1110111011100110",
    "1110100010110011",
    "1110001111101001",
    "1110000011011000",
    "1101111101110101",
    "1101111101010010",
    "1101111111001100",
    "1110000001010010",
    "1110000010110100",
    "1110000100100101",
    "1110001001011101",
    "1110010110011000",
    "1110101110111101",
    "1111010011000001",
    "1111111110001001",
    "1111010111100011",
    "1110110110010010",
    "1110100100000000",
    "1110100011000000",
    "1110110000001111",
    "1111000101010000",
    "1111011011101111",
    "1111101111111110",
    "1111111101101110",
    "1111101010110110",
    "1111010101011010",
    "1110111101001100",
    "1110100100010010",
    "1110001110110000",
    "1110000000011110",
    "1101111011110010",
    "1110000000011110",
    "1110001100000001",
    "1110011011011011",
    "1110101101100011",
    "1111000010111011",
    "1111011100001010",
    "1111111000000101",
    "1111101100101110",
    "1111010110110001",
    "1111001001111010",
    "1111001000010110",
    "1111010001010101",
    "1111100001111011",
    "1111110110010100",
    "1111110100111100",
    "1111100010011001",
    "1111010011011010",
    "1111001001010001",
    "1111000101100101",
    "1111001010011101",
    "1111011001101111",
    "1111110011100001",
    "1111101010101101",
    "1111000101111011",
    "1110100100001110",
    "1110001011011001",
    "1101111110101110",
    "1101111110010010",
    "1110000111010001",
    "1110010101111001",
    "1110100111100000",
    "1110111100000001",
    "1111010100111100",
    "1111110011011110",
    "1111101001011111",
    "1111000101101010",
    "1110100110000110",
    "1110001111101011",
    "1110000101001001",
    "1110000101101001",
    "1110001100111000",
    "1110010101101111",
    "1110011100001110",
    "1110011111000100",
    "1110011111100100",
    "1110100000010100",
    "1110100011101100",
    "1110101011101010",
    "1110111010000010",
    "1111010000000011",
    "1111101101001100",
    "1111110001001011",
    "1111001111110011",
    "1110110100001011",
    "1110100010110001",
    "1110011110000101",
    "1110100101000001",
    "1110110011000101",
    "1111000010010111",
    "1111001101110101",
    "1111010010110100",
    "1111010001100010",
    "1111001100001111",
    "1111000110001011",
    "1111000011100100",
    "1111001000101111",
    "1111011000000110",
    "1111110000111101",
    "1111110000101000",
    "1111010010110011",
    "1110111011011001",
    "1110101110110101",
    "1110101111000010",
    "1110111010011101",
    "1111001100101000",
    "1111011111111111",
    "1111101111100011",
    "1111111000100010",
    "1111111001111111",
    "1111110100001010",
    "1111101000011110",
    "1111011000110100",
    "1111000111001000",
    "1110110101110001",
    "1110100111001011",
    "1110011101100100",
    "1110011010101101",
    "1110011111000111",
    "1110101010101010",
    "1110111101011100",
    "1111010111100111",
    "1111111000011111",
    "1111100010011100",
    "1110111101110011",
    "1110011111000100",
    "1110001010101010",
    "1110000010111011",
    "1110000110101100",
    "1110010001110001",
    "1110011111001100",
    "1110101100000100",
    "1110111000111111",
    "1111001001000001",
    "1111011111000010",
    "1111111011110110",
    "1111100010101001",
    "1111000001000011",
    "1110100100101001",
    "1110010001011111",
    "1110001000110100",
    "1110001001010011",
    "1110010000001111",
    "1110011011000001",
    "1110101000001000",
    "1110110111001101",
    "1111000111101010",
    "1111011000000100",
    "1111100101110110",
    "1111101110001100",
    "1111101111010010",
    "1111101001000110",
    "1111011101011100",
    "1111001111011010",
    "1111000010011001",
    "1110111000110111",
    "1110110011111001",
    "1110110011000101",
    "1110110101100101",
    "1110111010111111",
    "1111000011111100",
    "1111010001111101",
    "1111100110001011",
    "1111111111011110",
    "1111100001000011",
    "1111000010000011",
    "1110100110100101",
    "1110010001101110",
    "1110000100101001",
    "1101111110111010",
    "1101111111000101",
    "1110000011101010",
    "1110001011100000",
    "1110010101110001",
    "1110100001101110",
    "1110101110011001",
    "1110111010100110",
    "1111000110000100",
    "1111010010110011",
    "1111100011101100",
    "1111111010011010",
    "1111101010011010",
    "1111001111101110",
    "1110111100000101",
    "1110110101110110",
    "1111000001001111",
    "1111011110000111",
    "1111111000011111",
    "1111001010011011",
    "1110100000000000",
    "1101111111101000",
    "1101101100010001",
    "1101100101110111",
    "1101101001111001",
    "1101110100011101",
    "1110000010101111",
    "1110010011111110",
    "1110101000110000",
    "1111000001110110",
    "1111011110010110",
    "1111111011000011",
    "1111101100001110",
    "1111011011001010",
    "1111010011001000",
    "1111010010100010",
    "1111010101100101",
    "1111010111110010",
    "1111010101110111",
    "1111001110111101",
    "1111000100110110",
    "1110111010100101",
    "1110110011010000",
    "1110110000011110",
    "1110110010000011",
    "1110110110100100",
    "1110111100010011",
    "1111000010101011",
    "1111001011010110",
    "1111011000111001",
    "1111101100100001",
    "1111111011001100",
    "1111100010110011",
    "1111001111100100",
    "1111000110000100",
    "1111001000100000",
    "1111010101101010",
    "1111101001001011",
    "1111111101011010",
    "1111110010111101",
    "1111101011010101",
    "1111101100011101",
    "1111110101010011",
    "1111111100000100",
    "1111101001110000",
    "1111010101001011",
    "1110111111100001",
    "1110101010000111",
    "1110010110100101",
    "1110000111000011",
    "1101111101011100",
    "1101111010111010",
    "1101111111000101",
    "1110001000001001",
    "1110010100000101",
    "1110100001001000",
    "1110101110011111",
    "1110111101100100",
    "1111010001110001",
    "1111101101100111",
    "1111101111000011",
    "1111001000001011",
    "1110100100010101",
    "1110001010010110",
    "1101111111000101",
    "1110000011110001",
    "1110010100110001",
    "1110101100000001",
    "1111000011100001",
    "1111010111010110",
    "1111100110011110",
    "1111110001011111",
    "1111111001001001",
    "1111111101110110",
    "1111111111000111",
    "1111111100000011",
    "1111110100100100",
    "1111101001100101",
    "1111011101000101",
    "1111010001111000",
    "1111001010101010",
    "1111001001000110",
    "1111001101101101",
    "1111010111111001",
    "1111100110100000",
    "1111110111110100",
    "1111110110011101",
    "1111100111000110",
    "1111011100101000",
    "1111011000101000",
    "1111011011001111",
    "1111100011010010",
    "1111101110111101",
    "1111111100000110",
    "1111110111001111",
    "1111101100100001",
    "1111100100001010",
    "1111011101101110",
    "1111011000110100",
    "1111010101000110",
    "1111010010110001",
    "1111010010100111",
    "1111010110000001",
    "1111011110001101",
    "1111101011101010",
    "1111111101010110",
    "1111101111000101",
    "1111011100100011",
    "1111001101100001",
    "1111000011100010",
    "1110111110101101",
    "1110111110000100",
    "1111000000001100",
    "1111000011100010",
    "1111000111010011",
    "1111001011000111",
    "1111001111001000",
    "1111010011010111",
    "1111010111101000",
    "1111011100000010",
    "1111100000111110",
    "1111100111000110",
    "1111101110111001",
    "1111111000010101",
    "1111111101001100",
    "1111110011001101",
    "1111101011110011",
    "1111101001010101",
    "1111101101101011",
    "1111111001011111",
    "1111110100011100",
    "1111011111001010",
    "1111001010101010",
    "1110111010110000",
    "1110110010010000",
    "1110110001111001",
    "1110111000010110",
    "1111000010110110",
    "1111001111000111",
    "1111011100101010",
    "1111101100001011",
    "1111111110001010",
    "1111101110001000",
    "1111011011011011",
    "1111001101011011",
    "1111000111110101",
    "1111001100111010",
    "1111011100000101",
    "1111110010001111",
    "1111110101010010",
    "1111011111010110",
    "1111001111010110",
    "1111000110111001",
    "1111000101110111",
    "1111001010100110",
    "1111010010011111",
    "1111011010101000",
    "1111100000010111",
    "1111100001101110",
    "1111011101111111",
    "1111010101101110",
    "1111001010100110",
    "1110111111000111",
    "1110110101110110",
    "1110110000110011",
    "1110110000111001",
    "1110110101101010",
    "1110111101110101",
    "1111001000100000",
    "1111010101101010",
    "1111100110000011",
    "1111111010000100",
    "1111101110111010",
    "1111010111000001",
    "1111000001010101",
    "1110110001001101",
    "1110101001000110",
    "1110101001011101",
    "1110110000101001",
    "1110111011100110",
    "1111000111000110",
    "1111010000110000",
    "1111011000011101",
    "1111100001001000",
    "1111101110100101",
    "1111111101000011",
    "1111100011000011",
    "1111000111111110",
    "1110110001110001",
    "1110100101100000",
    "1110100101010101",
    "1110101111011001",
    "1110111110110011",
    "1111001110001101",
    "1111011001100011",
    "1111011111011100",
    "1111100000101110",
    "1111011111010001",
    "1111011101000111",
    "1111011011100001",
    "1111011010100101",
    "1111011001110101",
    "1111011001001001",
    "1111011000111010",
    "1111011010011101",
    "1111011111100100",
    "1111101001011100",
    "1111110111110000",
    "1111110111001001",
    "1111100101101100",
    "1111010110000000",
    "1111001001101000",
    "1111000001001101",
    "1110111100011110",
    "1110111010100011",
    "1110111010011001",
    "1110111011000110",
    "1110111100000111",
    "1110111101010010",
    "1110111110101000",
    "1111000000001101",
    "1111000010010101",
    "1111000101100000",
    "1111001010001100",
    "1111010000110011",
    "1111011001011101",
    "1111100011110011",
    "1111101110110010",
    "1111111001010110",
    "1111111101010111",
    "1111110101101111",
    "1111101111101011",
    "1111101010111101",
    "1111100111011000",
    "1111100100111001",
    "1111100011100001",
    "1111100011000001",
    "1111100010111101",
    "1111100010110011",
    "1111100010101110",
    "1111100011101111",
    "1111100111101001",
    "1111110000000111",
    "1111111101111100",
    "1111101111110110",
    "1111011100001010",
    "1111001010111000",
    "1110111111110001",
    "1110111101010010",
    "1111000011101111",
    "1111010001001100",
    "1111100001111011",
    "1111110001011111",
    "1111111011110010",
    "1111111101110100",
    "1111110110010100",
    "1111100110000011",
    "1111001111101110",
    "1110110111010011",
    "1110100001001101",
    "1110010001000010",
    "1110001000101101",
    "1110001000001011",
    "1110001101010111",
    "1110010101101001",
    "1110011111111011",
    "1110101101011001",
    "1110111111101011",
    "1111010111001000",
    "1111110001100101",
    "1111110101010001",
    "1111100010010101",
    "1111011001010001",
    "1111011010111010",
    "1111100100011000",
    "1111110000111000",
    "1111111011101000",
    "1111111110000111",
    "1111111100011111",
    "1111111101101000",
    "1111111111000011",
    "1111111110011000",
    "1111111010011000",
    "1111110010110101",
    "1111100111111110",
    "1111011010011000",
    "1111001010110101",
    "1110111010011000",
    "1110101010101010",
    "1110011110001010",
    "1110010111100010",
    "1110011000111010",
    "1110100011001000",
    "1110110101101100",
    "1111001110110101",
    "1111101011011111",
    "1111111000000100",
    "1111011111110000",
    "1111001110110011",
    "1111000110111110",
    "1111001000000011",
    "1111001111111111",
    "1111011011011110",
    "1111100111000111",
    "1111110001001111",
    "1111111011010001",
    "1111110111100101",
    "1111100100111001",
    "1111001100100011",
    "1110110001110000",
    "1110011001101011",
    "1110001001110111",
    "1110000110001000",
    "1110001110100011",
    "1110011111011001",
    "1110110010110110",
    "1111000011011000",
    "1111001101101000",
    "1111010001000011",
    "1111001111000101",
    "1111001010001011",
    "1111000100101111",
    "1111000000001101",
    "1110111101010001",
    "1110111100000101",
    "1110111100010100",
    "1110111101010111",
    "1110111110110011",
    "1111000000010010",
    "1111000001101100",
    "1111000011000001",
    "1111000101000110",
    "1111001001100010",
    "1111010010010010",
    "1111100000100011",
    "1111110100000100",
    "1111110100111110",
    "1111011101110011",
    "1111001001111010",
    "1110111100000101",
    "1110110101011111",
    "1110110101001001",
    "1110111000101101",
    "1110111101011001",
    "1111000001000111",
    "1111000010111011",
    "1111000011000011",
    "1111000010001111",
    "1111000001001111",
    "1111000000101011",
    "1111000000101110",
    "1111000001100010",
    "1111000011011000",
    "1111000110011011",
    "1111001010100101",
    "1111001111001101",
    "1111010011010011",
    "1111010101110001",
    "1111010110000110",
    "1111010100101110",
    "1111010010111001",
    "1111010010010101",
    "1111010100011111",
    "1111011001111111",
    "1111100010010100",
    "1111101100000101",
    "1111110101110111",
    "1111111110110001",
    "1111111001001011",
    "1111110001101010",
    "1111101010011001",
    "1111100011011000",
    "1111011101000000",
    "1111011000000011",
    "1111010101001011",
    "1111010100101010",
    "1111010110010010",
    "1111011001100000",
    "1111011110011011",
    "1111100110000001",
    "1111110001111001",
    "1111111100111101",
    "1111100111010110",
    "1111001111111111",
    "1110111010101011",
    "1110101011001100",
    "1110100011111001",
    "1110100101000001",
    "1110101101010111",
    "1110111011011001",
    "1111001110000101",
    "1111100100100010",
    "1111111101010000",
    "1111101010011000",
    "1111010101110110",
    "1111001000011000",
    "1111000100010111",
    "1111001010100011",
    "1111011010011000",
    "1111110010001011",
    "1111110000100010",
    "1111010000111110",
    "1110110010011101",
    "1110011000001001",
    "1110000100101001",
    "1101111001111101",
    "1101111001101011",
    "1110000100110011",
    "1110011011011000",
    "1110111011101011",
    "1111100001101100",
    "1111111000000000",
    "1111010111001110",
    "1111000000000000",
    "1110110011110001",
    "1110110001000101",
    "1110110100011010",
    "1110111001110000",
    "1110111110000010",
    "1110111111110001",
    "1110111111010111",
    "1110111110010001",
    "1110111110010001",
    "1111000000101110",
    "1111000101100111",
    "1111001011110111",
    "1111010001110110",
    "1111010110000110",
    "1111011000100111",
    "1111011100010100",
    "1111100101000110",
    "1111110100111111",
    "1111110100110110",
    "1111011100011100",
    "1111000110111100",
    "1110111001000010",
    "1110110101110001",
    "1110111100101000",
    "1111001010010011",
    "1111011010110010",
    "1111101010110100",
    "1111111000100101",
    "1111111100010011",
    "1111110100000101",
    "1111101110111001",
    "1111101101000111",
    "1111101111110001",
    "1111110111101011",
    "1111111011001100",
    "1111101001101101",
    "1111010101011101",
    "1111000000011111",
    "1110101100110101",
    "1110011011111101",
    "1110001110111011",
    "1110000110101000",
    "1110000011100110",
    "1110000110000100",
    "1110001110100011",
    "1110011101101000",
    "1110110011010010",
    "1111001110000111",
    "1111101011010000",
    "1111111001010001",
    "1111100011011111",
    "1111010110010010",
    "1111010010101001",
    "1111010111100000",
    "1111100010101110",
    "1111110010000000",
    "1111111100011101",
    "1111101010000110",
    "1111011000001110",
    "1111001000110010",
    "1110111101111000",
    "1110111001010110",
    "1110111011111101",
    "1111000101000110",
    "1111010010111000",
    "1111100010111000",
    "1111110010100111",
    "1111111111011101",
    "1111110100000001",
    "1111101010110100",
    "1111100011001011",
    "1111011100110000",
    "1111010111110010",
    "1111010101000011",
    "1111010101100010",
    "1111011001111111",
    "1111100011000000",
    "1111110000101011",
    "1111111101011100",
    "1111101000100001",
    "1111010010000110",
    "1110111100000111",
    "1110101000100101",
    "1110011001100011",
    "1110010000111001",
    "1110010000000011",
    "1110010111110111",
    "1110101000011010",
    "1111000000011111",
    "1111011101011001",
    "1111111011001010",
    "1111101010010101",
    "1111010110101000",
    "1111001011110111",
    "1111001010011110",
    "1111010001101100",
    "1111011111101001",
    "1111110010010101",
    "1111111000011001",
    "1111100010101110",
    "1111001110100011",
    "1110111101110000",
    "1110110001111011",
    "1110101100001001",
    "1110101100110010",
    "1110110011101001",
    "1111000000101011",
    "1111010100010111",
    "1111101110111101",
    "1111110000100101",
    "1111001101010110",
    "1110101011110011",
    "1110010000111001",
    "1110000000110001",
    "1101111101101011",
    "1110001000000110",
    "1110011111010111",
    "1111000001111000",
    "1111101100011011",
    "1111100101100010",
    "1110111001101111",
    "1110010101110010",
    "1101111101111010",
    "1101110011111001",
    "1101110110010101",
    "1110000001010111",
    "1110010000010100",
    "1110011111010001",
    "1110101100111000",
    "1110111011001111",
    "1111001101100100",
    "1111100101111100",
    "1111111100010111",
    "1111011101111010",
    "1111000100110111",
    "1110110110111100",
    "1110110111010011",
    "1111000100100101",
    "1111011001100101",
    "1111101111101010",
    "1111111111000010",
    "1111110110000001",
    "1111110101111000",
    "1111111101011000",
    "1111110110010000",
    "1111101000010001",
    "1111011011001001",
    "1111010000100110",
    "1111001001011110",
    "1111000101111110",
    "1111000101110111",
    "1111001000101101",
    "1111001101011100",
    "1111010010011111",
    "1111010110001001",
    "1111010111011101",
    "1111010110011111",
    "1111010100001011",
    "1111010001111001",
    "1111010000111001",
    "1111010001111101",
    "1111010101010010",
    "1111011010101011",
    "1111100001100110",
    "1111101001001111",
    "1111110000110000",
    "1111110111011000",
    "1111111100100011",
    "1111111111110111",
    "1111111110000010",
    "1111111101110110",
    "1111111111010001",
    "1111111101110000",
    "1111111001100110",
    "1111110100100010",
    "1111101110101111",
    "1111101000000000",
    "1111100000000010",
    "1111010110100111",
    "1111001100000101",
    "1111000001010100",
    "1110110111011101",
    "1110110000000010",
    "1110101100011011",
    "1110101101110000",
    "1110110100111011",
    "1111000010001101",
    "1111010101001101",
    "1111101100100011",
    "1111111001111111",
    "1111100001001101",
    "1111001011110010",
    "1110111011101111",
    "1110110010000000",
    "1110101110010110",
    "1110101111100001",
    "1110110011110100",
    "1110111001100011",
    "1110111111010110",
    "1111000100010010",
    "1111001000000011",
    "1111001010011110",
    "1111001011101011",
    "1111001011110101",
    "1111001011011001",
    "1111001011000001",
    "1111001011100000",
    "1111001101100001",
    "1111010001010111",
    "1111010110110100",
    "1111011101010110",
    "1111100100100101",
    "1111101100100001",
    "1111110101100001",
    "1111111111110100",
    "1111110011001001",
    "1111100100011010",
    "1111010100001010",
    "1111000011001000",
    "1110110010001010",
    "1110100010000011",
    "1110010011101010",
    "1110000111111010",
    "1101111111110011",
    "1101111100010011",
    "1101111110000111",
    "1110000101100111",
    "1110010011000001",
    "1110100110100101",
    "1111000000000011",
    "1111011110100011",
    "1111111111110011",
    "1111011111101001",
    "1111000011101110",
    "1110101111101110",
    "1110100101011111",
    "1110100100101100",
    "1110101011000111",
    "1110110101100010",
    "1111000000110101",
    "1111001010110000",
    "1111010010100110",
    "1111011001011000",
    "1111100001111000",
    "1111101110110100",
    "1111111110101001",
    "1111101000001000",
    "1111010001100110",
    "1111000000010111",
    "1110111001011000",
    "1110111111011110",
    "1111010001111110",
    "1111101100110000",
    "1111110110001101",
    "1111011101000100",
    "1111001100001110",
    "1111000101011111",
    "1111001000001110",
    "1111010010001010",
    "1111100001001000",
    "1111110100001011",
    "1111110101000111",
    "1111011011100101",
    "1111000001010000",
    "1110101001110000",
    "1110011001001110",
    "1110010011000001",
    "1110011000010101",
    "1110100111011111",
    "1110111100110011",
    "1111010011100010",
    "1111100111000100",
    "1111110100000100",
    "1111111000110110",
    "1111110101011111",
    "1111101011101000",
    "1111011101110101",
    "1111001110111011",
    "1111000001100001",
    "1110110111011010",
    "1110110001110100",
    "1110110001100111",
    "1110110111011011",
    "1111000011000011",
    "1111010011010010",
    "1111100101101010",
    "1111110110111101",
    "1111111011111010",
    "1111110101010111",
    "1111110110010110",
    "1111111110011011",
    "1111110011101111",
    "1111100010000110",
    "1111001110110011",
    "1110111100000010",
    "1110101100001100",
    "1110100001011111",
    "1110011101010100",
    "1110011111111010",
    "1110100111111010",
    "1110110010101111",
    "1110111101100000",
    "1111000101110110",
    "1111001011000010",
    "1111001101111101",
    "1111010000010010",
    "1111010101000101",
    "1111100000110001",
    "1111110110011100",
    "1111101010010111",
    "1111000101111110",
    "1110100011010011",
    "1110001001010000",
    "1101111100101011",
    "1101111111010010",
    "1110001110001010",
    "1110100011010011",
    "1110111000100101",
    "1111001001001100",
    "1111010011010000",
    "1111010111001011",
    "1111010110100010",
    "1111010011100010",
    "1111010000000111",
    "1111001101000000",
    "1111001010100010",
    "1111001000101010",
    "1111000111100111",
    "1111001000101101",
    "1111001110010001",
    "1111011010000001",
    "1111101100000010",
    "1111111101101110",
    "1111100110110100",
    "1111010010111110",
    "1111000101011011",
    "1110111111111010",
    "1111000001101100",
    "1111001000010011",
    "1111010000011010",
    "1111010111011101",
    "1111011100100000",
    "1111100000010101",
    "1111100100101100",
    "1111101011010111",
    "1111110101011101",
    "1111111101010110",
    "1111101110100100",
    "1111100000011001",
    "1111010101000110",
    "1111001110100110",
    "1111001110010010",
    "1111010100111001",
    "1111100010001111",
    "1111110100111011",
    "1111110101010011",
    "1111011111010111",
    "1111001011110111",
    "1110111100110111",
    "1110110011101001",
    "1110110000101001",
    "1110110011101001",
    "1110111011110011",
    "1111000111110101",
    "1111010110100101",
    "1111100111000011",
    "1111111000011001",
    "1111110110001101",
    "1111100101100111",
    "1111010110101100",
    "1111001010010110",
    "1111000001100100",
    "1110111100101011",
    "1110111011011000",
    "1110111100110101",
    "1111000000001101",
    "1111000101001001",
    "1111001011011001",
    "1111010010011101",
    "1111011001010101",
    "1111011101111111",
    "1111011110000000",
    "1111010111001110",
    "1111001000111010",
    "1110110100100100",
    "1110011101110000",
    "1110001001000110",
    "1101111010101000",
    "1101110100100010",
    "1101110110100101",
    "1101111110101000",
    "1110001001101101",
    "1110010101011000",
    "1110100000100100",
    "1110101011110000",
    "1110111001111001",
    "1111001110111010",
    "1111101100110111",
    "1111101101011011",
    "1111000100110111",
    "1110100000001100",
    "1110000101011111",
    "1101111000100010",
    "1101111001011011",
    "1110000100010000",
    "1110010011010111",
    "1110100001110001",
    "1110101100100101",
    "1110110011011100",
    "1110110111011000",
    "1110111001111010",
    "1110111100010100",
    "1110111111001010",
    "1111000010000000",
    "1111000100101001",
    "1111001000111010",
    "1111010011001011",
    "1111100111001100",
    "1111111010010101",
    "1111010100111001",
    "1110101111011110",
    "1110010001011010",
    "1110000000001101",
    "1101111101100011",
    "1110000110010011",
    "1110010100101111",
    "1110100011101110",
    "1110110001100010",
    "1111000000011010",
    "1111010011100001",
    "1111101100010000",
    "1111110110101100",
    "1111011001110010",
    "1111000010100100",
    "1110110101011101",
    "1110110011111011",
    "1110111011110010",
    "1111001000110000",
    "1111010110110010",
    "1111100011101100",
    "1111101111100111",
    "1111111011010000",
    "1111111001101100",
    "1111110001000001",
    "1111101101010010",
    "1111110000100010",
    "1111111011000100",
    "1111110100110111",
    "1111100010110011",
    "1111010010101011",
    "1111000111100010",
    "1111000010011100",
    "1111000010010010",
    "1111000100111011",
    "1111001000101010",
    "1111001101100001",
    "1111010101101010",
    "1111100100000011",
    "1111111010001001",
    "1111101001010101",
    "1111001010111010",
    "1110110000101100",
    "1110100000010101",
    "1110011101000101",
    "1110100110101000",
    "1110111001101111",
    "1111010010000110",
    "1111101011111110",
    "1111111011000010",
    "1111100100001010",
    "1111001111110110",
    "1110111110100011",
    "1110110000110101",
    "1110100111100000",
    "1110100011001000",
    "1110100011010101",
    "1110100111010110",
    "1110101110101110",
    "1110111001100010",
    "1111001000011000",
    "1111011011111100",
    "1111110100000011",
    "1111110000110001",
    "1111010101010010",
    "1110111100101110",
    "1110101010000001",
    "1110011110100100",
    "1110011001111010",
    "1110011010001011",
    "1110011101000101",
    "1110100000110001",
    "1110100100011010",
    "1110101000000100",
    "1110101100100011",
    "1110110010100100",
    "1110111010000110",
    "1111000001111011",
    "1111001000001011",
    "1111001011000001",
    "1111001001011001",
    "1111000011011000",
    "1110111010010001",
    "1110110000001101",
    "1110100111101101",
    "1110100011000000",
    "1110100011110001",
    "1110101011001010",
    "1110111001110010",
    "1111001111101000",
    "1111101011100100",
    "1111110100110000",
    "1111010100110111",
    "1110111000101111",
    "1110100011111100",
    "1110011000111010",
    "1110011000000011",
    "1110011111011111",
    "1110101100000010",
    "1110111001111010",
    "1111000110110100",
    "1111010011100001",
    "1111100011001010",
    "1111111000101000",
    "1111101011010111",
    "1111001011100101",
    "1110101101000101",
    "1110010101011010",
    "1110001000110101",
    "1110001000010110",
    "1110010001000011",
    "1110011110000101",
    "1110101010101010",
    "1110110011110011",
    "1110111001000010",
    "1110111011011011",
    "1110111100101101",
    "1110111110100011",
    "1111000001110110",
    "1111000111000100",
    "1111001111001100",
    "1111011011100000",
    "1111101101001000",
    "1111111011110001",
    "1111100001001100",
    "1111000110110110",
    "1110110001010101",
    "1110100100100100",
    "1110100010001111",
    "1110101001111001",
    "1110111001100011",
    "1111001110001101",
    "1111100100010111",
    "1111111000101100",
    "1111110111011110",
    "1111101110000010",
    "1111101011110110",
    "1111110000110101",
    "1111111100010001",
    "1111110011001011",
    "1111011111100011",
    "1111001011000111",
    "1110111000010011",
    "1110101001001001",
    "1110011111001100",
    "1110011011000110",
    "1110011100101011",
    "1110100011101001",
    "1110110000011111",
    "1111000100011000",
    "1111011111100110",
    "1111111111100110",
    "1111011101010110",
    "1110111110101110",
    "1110101000011101",
    "1110011101010001",
    "1110011101010001",
    "1110100101110110",
    "1110110010110001",
    "1111000000011001",
    "1111001101100011",
    "1111011100001110",
    "1111101111010101",
    "1111110111011000",
    "1111011001001100",
    "1110111010010110",
    "1110100000100111",
    "1110010001101011",
    "1110010001000011",
    "1110011111001111",
    "1110111001100111",
    "1111011011100000",
    "1111111111100110",
    "1111011111000000",
    "1111000100011000",
    "1110110011010010",
    "1110101100111100",
    "1110110001001101",
    "1110111110110101",
    "1111010100000000",
    "1111101110011011",
    "1111110100100011",
    "1111011000000110",
    "1110111111010110",
    "1110101100110101",
    "1110100010001010",
    "1110011111110000",
    "1110100101001000",
    "1110110001001010",
    "1111000010001011",
    "1111010101111011",
    "1111101001111111",
    "1111111100010001",
    "1111110100101010",
    "1111101001011011",
    "1111100001111011",
    "1111011101101101",
    "1111011100010110",
    "1111011101101000",
    "1111100001110001",
    "1111101001101101",
    "1111110110101101",
    "1111110110010010",
    "1111011101110010",
    "1111000010000110",
    "1110100111010000",
    "1110010010000101",
    "1110000110101111",
    "1110000111100111",
    "1110010100101110",
    "1110101100001010",
    "1111001011000111",
    "1111101110000010",
    "1111101110101101",
    "1111001110101001",
    "1110110100110011",
    "1110100011001011",
    "1110011011000001",
    "1110011100001100",
    "1110100101011010",
    "1110110100001011",
    "1111000101010000",
    "1111010101100010",
    "1111100010011100",
    "1111101010110110",
    "1111110000001010",
    "1111110110011101",
    "1111111110000000",
    "1111101011001010",
    "1111010010011111",
    "1110111000101010",
    "1110100011110100",
    "1110011001100011",
    "1110011101001010",
    "1110101110001001",
    "1111001000101101",
    "1111100111010011",
    "1111111100000010",
    "1111100101111001",
    "1111011000111110",
    "1111010110100000",
    "1111011110010100",
    "1111101111011000",
    "1111111000001000",
    "1111011011000110",
    "1110111101000111",
    "1110100010010010",
    "1110001110011111",
    "1110000100011010",
    "1110000100011010",
    "1110001100011100",
    "1110011000111001",
    "1110100101110100",
    "1110110000000111",
    "1110110110000001",
    "1110110111000110",
    "1110110100001101",
    "1110101111000000",
    "1110101001010001",
    "1110100100101001",
    "1110100010001011",
    "1110100011101001",
    "1110101100000100",
    "1110111110000000",
    "1111011001011001",
    "1111111010101111",
    "1111100100010010",
    "1111001010100101",
    "1110111101011001",
    "1110111110100100",
    "1111001011001111",
    "1111011101001110",
    "1111101110000110",
    "1111111001101100",
    "1111111111101011",
    "1111111101010111",
    "1111111010010110",
    "1111110100111010",
    "1111101100101110",
    "1111100011100100",
    "1111011100000111",
    "1111011000101111",
    "1111011010101000",
    "1111100001010100",
    "1111101011010100",
    "1111110111100111",
    "1111111001111110",
    "1111101001011111",
    "1111010111011010",
    "1111000101001110",
    "1110110101000001",
    "1110101000111110",
    "1110100010111101",
    "1110100100001000",
    "1110101100100110",
    "1110111011011110",
    "1111001110110110",
    "1111100100001011",
    "1111111000101110",
    "1111110110001011",
    "1111101010111010",
    "1111100111000111",
    "1111101011011001",
    "1111110110110011",
    "1111111001000100",
    "1111100111111100",
    "1111011001111100",
    "1111010010101011",
    "1111010100001010",
    "1111011110001001",
    "1111101110010001",
    "1111111110111111",
    "1111101101010001",
    "1111011111001111",
    "1111010110000110",
    "1111010001101100",
    "1111010000101011",
    "1111010001010111",
    "1111010010010111",
    "1111010011001101",
    "1111010100001000",
    "1111010101101110",
    "1111011000010001",
    "1111011011111000",
    "1111100000010100",
    "1111100101000110",
    "1111101001100111",
    "1111101101001111",
    "1111101111100000",
    "1111110000010000",
    "1111101111011001",
    "1111101101000100",
    "1111101001100011",
    "1111100101001110",
    "1111100000100001",
    "1111011011110101",
    "1111010111100101",
    "1111010100000110",
    "1111010001101110",
    "1111010000100110",
    "1111010000110101",
    "1111010010100001",
    "1111010110000000",
    "1111011100001100",
    "1111100110001101",
    "1111110100100100",
    "1111111001000101",
    "1111100100100111",
    "1111010000100111",
    "1111000000000010",
    "1110110101001101",
    "1110110001000011",
    "1110110010110011",
    "1110111000100000",
    "1110111111111010",
    "1111000111100010",
    "1111001111010110",
    "1111011000010110",
    "1111100011110110",
    "1111110010010010",
    "1111111101011111",
    "1111101110000111",
    "1111100010101100",
    "1111011101111011",
    "1111100001001111",
    "1111101100110001",
    "1111111111110101",
    "1111100111000001",
    "1111001001110101",
    "1110101011000100",
    "1110001101110011",
    "1101110101011011",
    "1101100100110110",
    "1101011101101000",
    "1101011111100011",
    "1101101000100011",
    "1101110110110100",
    "1110001001101111",
    "1110100001100001",
    "1110111110000100",
    "1111011101100011",
    "1111111100011100",
    "1111101001100111",
    "1111011000100111",
    "1111010010100110",
    "1111010110010011",
    "1111011111111101",
    "1111101010111111",
    "1111110011100001",
    "1111110111111111",
    "1111111000111001",
    "1111110111111001",
    "1111110110111011",
    "1111110111010001",
    "1111111000111100",
    "1111111011011111",
    "1111111111010110",
    "1111111001010101",
    "1111101100001010",
    "1111011000010000",
    "1110111111101000",
    "1110100110111011",
    "1110010011100110",
    "1110001001111100",
    "1110001011010100",
    "1110010101010101",
    "1110100011001011",
    "1110101111110000",
    "1110110111010101",
    "1110111000101100",
    "1110110100101001",
    "1110101101000100",
    "1110100100101001",
    "1110011110010010",
    "1110011100110011",
    "1110100001111110",
    "1110101101111111",
    "1110111111010001",
    "1111010010110110",
    "1111100101010011",
    "1111110011001101",
    "1111111010001101",
    "1111111001111101",
    "1111110100010101",
    "1111101100100010",
    "1111100101110111",
    "1111100010011101",
    "1111100011001011",
    "1111100111101011",
    "1111101110110011",
    "1111110111011001",
    "1111111111100010",
    "1111110110110101",
    "1111101111000101",
    "1111101001000000",
    "1111100101100101",
    "1111100110000000",
    "1111101010111011",
    "1111110100000011",
    "1111111111111000",
    "1111110011111001",
    "1111101001111100",
    "1111100100001110",
    "1111100011011100",
    "1111100110110010",
    "1111101100010101",
    "1111110001110001",
    "1111110101001111",
    "1111110101101100",
    "1111110010110011",
    "1111101100110011",
    "1111100100011010",
    "1111011010110101",
    "1111010001100100",
    "1111001010000110",
    "1111000101101100",
    "1111000101000110",
    "1111001000011000",
    "1111001110011111",
    "1111010101100111",
    "1111011011101000",
    "1111011110111111",
    "1111011111000000",
    "1111011100000010",
    "1111010111001001",
    "1111010010000010",
    "1111001110100110",
    "1111001110100100",
    "1111010011001000",
    "1111011100100110",
    "1111101010010010",
    "1111111010100011",
    "1111110100110110",
    "1111100110001101",
    "1111011010111100",
    "1111010011010101",
    "1111001110011011",
    "1111001010101011",
    "1111000110100010",
    "1111000001000010",
    "1110111010000100",
    "1110110010011010",
    "1110101011000111",
    "1110100101000110",
    "1110100000110110",
    "1110011110100100",
    "1110011110111111",
    "1110100011001000",
    "1110101011110101",
    "1110111000111001",
    "1111001000010101",
    "1111010110100101",
    "1111011111100100",
    "1111100000000111",
    "1111010111010000",
    "1111000111000011",
    "1110110011111110",
    "1110100011010111",
    "1110011010000100",
    "1110011011000010",
    "1110100111000001",
    "1110111100010001",
    "1111010111001011",
    "1111110011001100",
    "1111110011111110",
    "1111100001100110",
    "1111010111001011",
    "1111010100011100",
    "1111010111111010",
    "1111011111100110",
    "1111101001011110",
    "1111110100010001",
    "1111111111100011",
    "1111110100101010",
    "1111101000011100",
    "1111011100001110",
    "1111010000111011",
    "1111000111101010",
    "1111000001001000",
    "1110111101001001",
    "1110111010100101",
    "1110110111101101",
    "1110110010111110",
    "1110101011101111",
    "1110100010100100",
    "1110011001001100",
    "1110010001110100",
    "1110001110011111",
    "1110010000011111",
    "1110011000101000",
    "1110100111101111",
    "1110111101111011",
    "1111011010000100",
    "1111111001001010",
    "1111101001001011",
    "1111010001100100",
    "1111000011011100",
    "1111000000000011",
    "1111000101110001",
    "1111010000100011",
    "1111011011101111",
    "1111100011101100",
    "1111100111011110",
    "1111101001001100",
    "1111101100111011",
    "1111110110100100",
    "1111111000001100",
    "1111100001000000",
    "1111000111111110",
    "1110110010001111",
    "1110100100000000",
    "1110011111000000",
    "1110100010000010",
    "1110101010001001",
    "1110110100000000",
    "1110111101001110",
    "1111000101011000",
    "1111001110000000",
    "1111011001101000",
    "1111101001111011",
    "1111111110100110",
    "1111101010110110",
    "1111010110011010",
    "1111000111111100",
    "1111000001111000",
    "1111000011111001",
    "1111001011100000",
    "1111010100111011",
    "1111011100100110",
    "1111011111111011",
    "1111011101110011",
    "1111010110100000",
    "1111001011101010",
    "1110111111110110",
    "1110110101101110",
    "1110101111001100",
    "1110101101000100",
    "1110101110101001",
    "1110110010011111",
    "1110110110111110",
    "1110111010110111",
    "1110111101110000",
    "1111000000110101",
    "1111000110111110",
    "1111010011100010",
    "1111101000011000",
    "1111111011000001",
    "1111011010000100",
    "1110111001101101",
    "1110011110110001",
    "1110001100100000",
    "1110000011010011",
    "1110000001101100",
    "1110000101010101",
    "1110001100010100",
    "1110010110001001",
    "1110100011010010",
    "1110110100010010",
    "1111001000111111",
    "1111011111110101",
    "1111110101111011",
    "1111111000001010",
    "1111101101100100",
    "1111101011111001",
    "1111110010110010",
    "1111111111101100",
    "1111101110011100",
    "1111011100001001",
    "1111001011001010",
    "1110111101010100",
    "1110110100000001",
    "1110110000001100",
    "1110110001110100",
    "1110111000001000",
    "1111000001100001",
    "1111001100110000",
    "1111011010001001",
    "1111101011000110",
    "1111111111010101",
    "1111100101110010",
    "1111001011001110",
    "1110110100001010",
    "1110100101010111",
    "1110100010011010",
    "1110101100101101",
    "1111000011001011",
    "1111100011000101",
    "1111110111101011",
    "1111010001110011",
    "1110101111110011",
    "1110010101110110",
    "1110000110110100",
    "1110000011101010",
    "1110001011011001",
    "1110011011000001",
    "1110101110111011",
    "1111000101101110",
    "1111100000010101",
    "1111111111101010",
    "1111011010011001",
    "1110110010011101",
    "1110001100110111",
    "1101101111100001",
    "1101011111111010",
    "1101100000001101",
    "1101101101111011",
    "1110000011100100",
    "1110011010111111",
    "1110110000000101",
    "1111000010010010",
    "1111010011011000",
    "1111100101100010",
    "1111111001111100",
    "1111110000010100",
    "1111011100001001",
    "1111001100011100",
    "1111000011010111",
    "1111000000111001",
    "1111000011010010",
    "1111001000000011",
    "1111001101011001",
    "1111010011001010",
    "1111011010011101",
    "1111100100100101",
    "1111110010001111",
    "1111111101010000",
    "1111101100000100",
    "1111011100111101",
    "1111010010001011",
    "1111001100110000",
    "1111001011111101",
    "1111001110000010",
    "1111010001010010",
    "1111010100111100",
    "1111011001000100",
    "1111011110000010",
    "1111100100000000",
    "1111101010010001",
    "1111101111100100",
    "1111110010010011",
    "1111110001011010",
    "1111101100110100",
    "1111100101001110",
    "1111011011110101",
    "1111010001110000",
    "1111001000001001",
    "1111000000000101",
    "1110111010100110",
    "1110111000100010",
    "1110111010010011",
    "1110111111110001",
    "1111001000011010",
    "1111010011011111",
    "1111100000100011",
    "1111101111011000",
    "1111111111111000",
    "1111101101011001",
    "1111011001110000",
    "1111000110100000",
    "1110110101100111",
    "1110101001000110",
    "1110100010010000",
    "1110100001011001",
    "1110100101110010",
    "1110101110101001",
    "1110111100001010",
    "1111001111010010",
    "1111101000101001",
    "1111111000100111",
    "1111010111011101",
    "1110110111111110",
    "1110011110100001",
    "1110001110100100",
    "1110001001010001",
    "1110001101010111",
    "1110011000001001",
    "1110100110100000",
    "1110110110001110",
    "1111000110000011",
    "1111010101011010",
    "1111100011111110",
    "1111110001011011",
    "1111111101010000",
    "1111111001000000",
    "1111110001110101",
    "1111101101011100",
    "1111101011101011",
    "1111101011111110",
    "1111101101101101",
    "1111110000010100",
    "1111110011010101",
    "1111110101111000",
    "1111110110011011",
    "1111110011001010",
    "1111101010110100",
    "1111011101000101",
    "1111001011001001",
    "1110110111001001",
    "1110100011111100",
    "1110010100001000",
    "1110001001100011",
    "1110000100111110",
    "1110000110010010",
    "1110001100110010",
    "1110010111101101",
    "1110100110010011",
    "1110111000001000",
    "1111001101011100",
    "1111100110110101",
    "1111111011100110",
    "1111011011001111",
    "1110111010111101",
    "1110011110011100",
    "1110001001001100",
    "1101111101100011",
    "1101111011111111",
    "1110000011001101",
    "1110010001010000",
    "1110100100110111",
    "1110111101100110",
    "1111011011000100",
    "1111111011110010",
    "1111100011001000",
    "1111000101101100",
    "1110101111101011",
    "1110100011011111",
    "1110100001011111",
    "1110101000100101",
    "1110110111100011",
    "1111001101011001",
    "1111101000111100",
    "1111110111110010",
    "1111011000010000",
    "1110111100110010",
    "1110101001111111",
    "1110100011101010",
    "1110101011101000",
    "1111000001000000",
    "1111100000001000",
    "1111111100100011",
    "1111011011010110",
    "1111000001011110",
    "1110110010000011",
    "1110101101100110",
    "1110110010001111",
    "1110111100101101",
    "1111001001100111",
    "1111010110001000",
    "1111100000101100",
    "1111101000110011",
    "1111101110110001",
    "1111110011111101",
    "1111111010101001",
    "1111111011000011",
    "1111101100100000",
    "1111011010101111",
    "1111001000100000",
    "1110111001010001",
    "1110110000000101",
    "1110101110100100",
    "1110110100011101",
    "1110111111110000",
    "1111001101101000",
    "1111011011100000",
    "1111100111111100",
    "1111110011010010",
    "1111111111000100",
    "1111110011001101",
    "1111100011010101",
    "1111010010110011",
    "1111000100010010",
    "1110111010100101",
    "1110110111010110",
    "1110111010100101",
    "1111000010100110",
    "1111001100111111",
    "1111010111110001",
    "1111100001111110",
    "1111101011111000",
    "1111110110110000",
    "1111111011101101",
    "1111101010001111",
    "1111010100101110",
    "1110111100101000",
    "1110100100110111",
    "1110010000101100",
    "1110000010111101",
    "1101111101000111",
    "1101111111010111",
    "1110001000111010",
    "1110011000100011",
    "1110101100111111",
    "1111000100110011",
    "1111011110001100",
    "1111110110110001",
    "1111110100001110",
    "1111100101011011",
    "1111011110100001",
    "1111011111111000",
    "1111101000011110",
    "1111110110000100",
    "1111111010000111",
    "1111101010110111",
    "1111011110001010",
    "1111010101010011",
    "1111010000110101",
    "1111010000111011",
    "1111010101011101",
    "1111011101111011",
    "1111101001011110",
    "1111110110110000",
    "1111111011100001",
    "1111101110101000",
    "1111100011101010",
    "1111011011110000",
    "1111011000001100",
    "1111011010100011",
    "1111100100000001",
    "1111110100110000",
    "1111110100100111",
    "1111011010110101",
    "1111000001010100",
    "1110101011000111",
    "1110011010010110",
    "1110001111101000",
    "1110001010001110",
    "1110001000110100",
    "1110001010001100",
    "1110001101101101",
    "1110010011010000",
    "1110011011011001",
    "1110100111100010",
    "1110111001100010",
    "1111010010010111",
    "1111110001000001",
    "1111101101110010",
    "1111001110111101",
    "1110110111011011",
    "1110101010110111",
    "1110101010100011",
    "1110110100101110",
    "1111000101100000",
    "1111011000101101",
    "1111101010110111",
    "1111111010010011",
    "1111111001010100",
    "1111101111111000",
    "1111101001001100",
    "1111100101101010",
    "1111100110010101",
    "1111101100100000",
    "1111111000111100",
    "1111110100101001",
    "1111011110010001",
    "1111000111000001",
    "1110110010011001",
    "1110100011010011",
    "1110011011101011",
    "1110011100110010",
    "1110100111111001",
    "1110111101111111",
    "1111011110011011",
    "1111111001110111",
    "1111010000001111",
    "1110101011001010",
    "1110010000011110",
    "1110000011101010",
    "1110000100110111",
    "1110010000100111",
    "1110100001110001",
    "1110110011011111",
    "1111000010110011",
    "1111001110111010",
    "1111011000100101",
    "1111100001001010",
    "1111101010000101",
    "1111110101000111",
    "1111111011111011",
    "1111101000101011",
    "1111010010001111",
    "1110111011100001",
    "1110101000001100",
    "1110011011011011",
    "1110010111001110",
    "1110011011100001",
    "1110100101101001",
    "1110110001011110",
    "1110111011001111",
    "1111000000101011",
    "1111000001011110",
    "1110111110011011",
    "1110111001000010",
    "1110110010111110",
    "1110101101010001",
    "1110101001000100",
    "1110101001010000",
    "1110110001010000",
    "1111000010111011",
    "1111011101001110",
    "1111111011011101",
    "1111101000111000",
    "1111010110000001",
    "1111001111110011",
    "1111010101111001",
    "1111100100000101",
    "1111110101001111",
    "1111111010100011",
    "1111101100110110",
    "1111100000101011",
    "1111010100100101",
    "1111000111111110",
    "1110111011100101",
    "1110110001101011",
    "1110101100111010",
    "1110101110110110",
    "1110110111101101",
    "1111000110001000",
    "1111010111111100",
    "1111101010101100",
    "1111111100100011",
    "1111110011011010",
    "1111100101100101",
    "1111011010001110",
    "1111010001011110",
    "1111001011001111",
    "1111000111001011",
    "1111000100100100",
    "1111000010110001",
    "1111000001101001",
    "1111000001010111",
    "1111000010001011",
    "1111000100010011",
    "1111000111100000",
    "1111001011000001",
    "1111001101100110",
    "1111001101111101",
    "1111001011010001",
    "1111000101100100",
    "1110111101110010",
    "1110110101110010",
    "1110110000001000",
    "1110110000000010",
    "1110111000110010",
    "1111001100011011",
    "1111101010101000",
    "1111101111100111",
    "1111000111011111",
    "1110100010100111",
    "1110000101111110",
    "1101110100001011",
    "1101101101000111",
    "1101101110100001",
    "1101110101001000",
    "1101111101110101",
    "1110000110100101",
    "1110001110000101",
    "1110010011110110",
    "1110011000001000",
    "1110011011001110",
    "1110011101100011",
    "1110011111011010",
    "1110100001000101",
    "1110100010111000",
    "1110100101000011",
    "1110100111100011",
    "1110101001111101",
    "1110101011101010",
    "1110101100001110",
    "1110101011111010",
    "1110101011100101",
    "1110101100001110",
    "1110101110101001",
    "1110110011010000",
    "1110111010101111",
    "1111000110100101",
    "1111011000011011",
    "1111110000100111",
    "1111110010010101",
    "1111010100001101",
    "1110111001101101",
    "1110100111010000",
    "1110011111101110",
    "1110100011001101",
    "1110101111001100",
    "1110111111110001",
    "1111010000110110",
    "1111011111100001",
    "1111101010100011",
    "1111110011010010",
    "1111111101001000",
    "1111110100110011",
    "1111100001111001",
    "1111001100100101",
    "1110111001101101",
    "1110101110110101",
    "1110110000000111",
    "1110111111001010",
    "1111011010000100",
    "1111111100011000",
    "1111011111010111",
    "1110111110011111",
    "1110100100100100",
    "1110010011001111",
    "1110001010011110",
    "1110001000111001",
    "1110001100100110",
    "1110010100000101",
    "1110011110010110",
    "1110101010111111",
    "1110111001111010",
    "1111001010111010",
    "1111011101011100",
    "1111110000110010",
    "1111111011111101",
    "1111101001111111",
    "1111011010100011",
    "1111001110101000",
    "1111000110100101",
    "1111000010000010",
    "1111000000001000",
    "1111000000000011",
    "1111000001010000",
    "1111000011010010",
    "1111000101110010",
    "1111001000011000",
    "1111001010101101",
    "1111001100100000",
    "1111001101111010",
    "1111010001001000",
    "1111011010001011",
    "1111101011111101",
    "1111111001011111",
    "1111011010000010",
    "1110111100001100",
    "1110100110101010",
    "1110011110101001",
    "1110100101110111",
    "1110111001101000",
    "1111010100100000",
    "1111110000011111",
    "1111110111011011",
    "1111100110000000",
    "1111011011110011",
    "1111011000001011",
    "1111011001010110",
    "1111011101101101",
    "1111100100001011",
    "1111101100010111",
    "1111110111000010",
    "1111111010101010",
    "1111101000100011",
    "1111010011110100",
    "1110111111000000",
    "1110101101010111",
    "1110100010001111",
    "1110100000011110",
    "1110101001100000",
    "1110111100110010",
    "1111010111110010",
    "1111110110111000",
    "1111101001111010",
    "1111001110000010",
    "1110110111111010",
    "1110101001000010",
    "1110100001101001",
    "1110100001000000",
    "1110100101101111",
    "1110101111000000",
    "1110111101010111",
    "1111010001111000",
    "1111101100111100",
    "1111110010101111",
    "1111010000111101",
    "1110110010110011",
    "1110011101100001",
    "1110010100101010",
    "1110011000110101",
    "1110100111110001",
    "1110111101101000",
    "1111010110010011",
    "1111101110100001",
    "1111111100000011",
    "1111101011010011",
    "1111100000101011",
    "1111011101011100",
    "1111100010100001",
    "1111101111111101",
    "1111111011011110",
    "1111100010100001",
    "1111001000110101",
    "1110110010001011",
    "1110100001001111",
    "1110010111001000",
    "1110010011010111",
    "1110010100011100",
    "1110011000110101",
    "1110100000000011",
    "1110101011000110",
    "1110111011011000",
    "1111010001100100",
    "1111101100100100",
    "1111110110101010",
    "1111011100101000",
    "1111001001011011",
    "1110111111101000",
    "1110111111001100",
    "1111000110001000",
    "1111010001010010",
    "1111011101110101",
    "1111101001111010",
    "1111110100111010",
    "1111111111100011",
    "1111110011111010",
    "1111100011010000",
    "1111001101111000",
    "1110110101101100",
    "1110011110110101",
    "1110001110001101",
    "1110000111101111",
    "1110001101000100",
    "1110011100100110",
    "1110110001111001",
    "1111000111011111",
    "1111011001001001",
    "1111100110000100",
    "1111110000010100",
    "1111111010101001",
    "1111111001010011",
    "1111101100010001",
    "1111100001010101",
    "1111011100100101",
    "1111100001011001",
    "1111110000100111",
    "1111111000001110",
    "1111011110001010",
    "1111000110101100",
    "1110110101111001",
    "1110101101101001",
    "1110101110000100",
    "1110110110000000",
    "1111000011100100",
    "1111010100101111",
    "1111100111101000",
    "1111111010100010",
    "1111110011110010",
    "1111100100100000",
    "1111011000100010",
    "1111010000010100",
    "1111001011100011",
    "1111001001001110",
    "1111001000000100",
    "1111000110111100",
    "1111000101001110",
    "1111000010110011",
    "1111000000001100",
    "1110111110100011",
    "1110111111110000",
    "1111000101111110",
    "1111010010110110",
    "1111100110011011",
    "1111111110110100",
    "1111100111011011",
    "1111010000110001",
    "1111000001000010",
    "1110111010011011",
    "1110111100101011",
    "1111000101001011",
    "1111010000001101",
    "1111011010010001",
    "1111100001000011",
    "1111100100100101",
    "1111100111011100",
    "1111101101000111",
    "1111111000000001",
    "1111111000001001",
    "1111100110101001",
    "1111011000010000",
    "1111010001101001",
    "1111010101110010",
    "1111100100100100",
    "1111111010111111",
    "1111101011101000",
    "1111010100000110",
    "1111000001111001",
    "1110110110100111",
    "1110110010011001",
    "1110110100011101",
    "1110111100010011",
    "1111001001111010",
    "1111011101100100",
    "1111110110111000",
    "1111101011101110",
    "1111001101100001",
    "1110110010110001",
    "1110011111010111",
    "1110010101101010",
    "1110010101101100",
    "1110011101010001",
    "1110101001001001",
    "1110110101111110",
    "1111000010111000",
    "1111010010000011",
    "1111100110011100",
    "1111111110110100",
    "1111011111110110",
    "1111000010000000",
    "1110101011100000",
    "1110100001011110",
    "1110100101110110",
    "1110110101111110",
    "1111001100110101",
    "1111100101110010",
    "1111111101111110",
    "1111101011001001",
    "1111010101010011",
    "1111000000101011",
    "1110101110001101",
    "1110011111110001",
    "1110010111100000",
    "1110010110100111",
    "1110011101000100",
    "1110101001110100",
    "1110111010111000",
    "1111001110001111",
    "1111100010010010",
    "1111110101110000",
    "1111111000101101",
    "1111101011010010",
    "1111100100010011",
    "1111100101011010",
    "1111101110110000",
    "1111111111000101",
    "1111101100001001",
    "1111010101111110",
    "1111000001000101",
    "1110101111011001",
    "1110100001110110",
    "1110011000101100",
    "1110010011110011",
    "1110010011000101",
    "1110010110011101",
    "1110011101101001",
    "1110101000000110",
    "1110110100111100",
    "1111000011010101",
    "1111010011010101",
    "1111100110001110",
    "1111111101100100",
    "1111100110011110",
    "1111001000010000",
    "1110101100001010",
    "1110010111100000",
    "1110001110011110",
    "1110010010011001",
    "1110100001000000",
    "1110110101111110",
    "1111001101001111",
    "1111100100011000",
    "1111111010110000",
    "1111101111101001",
    "1111011011100101",
    "1111001010111010",
    "1111000000111011",
    "1111000001101110",
    "1111001111110011",
    "1111101010100100",
    "1111110001111011",
    "1111001100010100",
    "1110101011100101",
    "1110010101000000",
    "1110001010101111",
    "1110001011011001",
    "1110010011010111",
    "1110011110011011",
    "1110101001000110",
    "1110110001011100",
    "1110111000000001",
    "1110111111111011",
    "1111001100111100",
    "1111100001011010",
    "1111111100101100",
    "1111100100110111",
    "1111001000110100",
    "1110110100010011",
    "1110101010100000",
    "1110101011000010",
    "1110110010101001",
    "1110111100111010",
    "1111000110010011",
    "1111001101011110",
    "1111010011011111",
    "1111011010110111",
    "1111100110010011",
    "1111110111000100",
    "1111110100010111",
    "1111011111111011",
    "1111010000010100",
    "1111001001010101",
    "1111001100001100",
    "1111010111001101",
    "1111100110110110",
    "1111110111100000",
    "1111111001001100",
    "1111101100001101",
    "1111100001011111",
    "1111011000100011",
    "1111010001010000",
    "1111001100001100",
    "1111001010100110",
    "1111001101110111",
    "1111010110110100",
    "1111100101001101",
    "1111110111101101",
    "1111110011100111",
    "1111011111001000",
    "1111001100110101",
    "1110111110001001",
    "1110110011111001",
    "1110101110011001",
    "1110101101101001",
    "1110110001011010",
    "1110111001000100",
    "1111000011111000",
    "1111010001010100",
    "1111100001000010",
    "1111110010110001",
    "1111111001111111",
    "1111100110011110",
    "1111010100011111",
    "1111000110000110",
    "1110111100111101",
    "1110111001110100",
    "1110111100001111",
    "1111000010110100",
    "1111001011011001",
    "1111010011100100",
    "1111011001011110",
    "1111011100001100",
    "1111011011011000",
    "1111010111000110",
    "1111001111100001",
    "1111000101000110",
    "1110111000101101",
    "1110101011101011",
    "1110011111100011",
    "1110010101110110",
    "1110001111101100",
    "1110001101011100",
    "1110001110011100",
    "1110010001100110",
    "1110010101101111",
    "1110011010011001",
    "1110100000101100",
    "1110101011001010",
    "1110111100000101",
    "1111010100001000",
    "1111110001010111",
    "1111110000010110",
    "1111010110010010",
    "1111000100110111",
    "1110111110011001",
    "1111000001111110",
    "1111001100011011",
    "1111011001110000",
    "1111100110101011",
    "1111110001001000",
    "1111111000011110",
    "1111111100111110",
    "1111111111001111",
    "1111111111100011",
    "1111111101101001",
    "1111111000111011",
    "1111110001001000",
    "1111100110101000",
    "1111011010101101",
    "1111001111000111",
    "1111000101100000",
    "1110111110110101",
    "1110111011001001",
    "1110111001110101",
    "1110111001110010",
    "1110111001101011",
    "1110111000100011",
    "1110110110000011",
    "1110110010101100",
    "1110101111101011",
    "1110101110101110",
    "1110110001110001",
    "1110111010100110",
    "1111001010000111",
    "1111011111101001",
    "1111111000110100",
    "1111101110001010",
    "1111011001100011",
    "1111001100110101",
    "1111001010000001",
    "1111010001010100",
    "1111100001101100",
    "1111111001001000",
    "1111101011001001",
    "1111001110101000",
    "1110110101000000",
    "1110100001110110",
    "1110010111101111",
    "1110010111100101",
    "1110100000001101",
    "1110101110111000",
    "1111000001100110",
    "1111011000000110",
    "1111110010110000",
    "1111101110101110",
    "1111001110011011",
    "1110101111111011",
    "1110010111010101",
    "1110001000010001",
    "1110000100011111",
    "1110001010100010",
    "1110010110110010",
    "1110100101000001",
    "1110110001111110",
    "1110111100011011",
    "1111000100110001",
    "1111001100001001",
    "1111010011111011",
    "1111011101101011",
    "1111101011010111",
    "1111111110011100",
    "1111101001010011",
    "1111001110010100",
    "1110110100101100",
    "1110100000111001",
    "1110010110110111",
    "1110011000011010",
    "1110100100000000",
    "1110110101010010",
    "1111000110110001",
    "1111010100000000",
    "1111011010111111",
    "1111011100000101",
    "1111011001000110",
    "1111010101000110",
    "1111010100100010",
    "1111011011101101",
    "1111101100100111",
    "1111111010000000",
    "1111011100100011",
    "1111000000100111",
    "1110101011001110",
    "1110011111101011",
    "1110011110011001",
    "1110100100100100",
    "1110101101111011",
    "1110110110101100",
    "1110111101011001",
    "1111000011100010",
    "1111001011110011",
    "1111011000010101",
    "1111101001001111",
    "1111111100000011",
    "1111110011011100",
    "1111101001101111",
    "1111101001110111",
    "1111110011101110",
    "1111111100000001",
    "1111101010011111",
    "1111011100001110",
    "1111010011111011",
    "1111010010001000",
    "1111010101101010",
    "1111011011111111",
    "1111100010100001",
    "1111100111110011",
    "1111101100000011",
    "1111110000101101",
    "1111110111001101",
    "1111111111111101",
    "1111110101110011",
    "1111101011110000",
    "1111100011101110",
    "1111011111010100",
    "1111011111101110",
    "1111100101011011",
    "1111110000010010",
    "1111111111011101",
    "1111101110001001",
    "1111011010001011",
    "1111000110101100",
    "1110110101110110",
    "1110101001011110",
    "1110100010101110",
    "1110100010001010",
    "1110100111111110",
    "1110110100000001",
    "1111000101101010",
    "1111011011100011",
    "1111110011101110",
    "1111110100000100",
    "1111011110001001",
    "1111001100001010",
    "1110111111001111",
    "1110110111001011",
    "1110110010110100",
    "1110110000011111",
    "1110101111000010",
    "1110101110001001",
    "1110101110011100",
    "1110110001000101",
    "1110110111001011",
    "1111000001010100",
    "1111001110111101",
    "1111011110010111",
    "1111101100111101",
    "1111111000001011",
    "1111111110000010",
    "1111111101011011",
    "1111110110011011",
    "1111101010010110",
    "1111011011100011",
    "1111001101000111",
    "1111000010010010",
    "1110111101110010",
    "1111000001110000",
    "1111001111001100",
    "1111100101100111",
    "1111111101010110",
    "1111011101111010",
    "1111000000110110",
    "1110101010101011",
    "1110011110010110",
    "1110011100101110",
    "1110100101000011",
    "1110110110010110",
    "1111010000011010",
    "1111110010111011",
    "1111100011110011",
    "1110110111100011",
    "1110001101110111",
    "1101101100100001",
    "1101011000001000",
    "1101010010001011",
    "1101011000100101",
    "1101100110101111",
    "1101110111100101",
    "1110000111000110",
    "1110010011011100",
    "1110011100100110",
    "1110100011110001",
    "1110101011000001",
    "1110110101000001",
    "1111000100000110",
    "1111011000111110",
    "1111110010010111",
    "1111110010110101",
    "1111011010110010",
    "1111001001010001",
    "1111000001000010",
    "1111000010011010",
    "1111001011000010",
    "1111010110110010",
    "1111100001000011",
    "1111100110100001",
    "1111100101111100",
    "1111011111111000",
    "1111010111011010",
    "1111010010001000",
    "1111010101100010",
    "1111100100011101",
    "1111111101110101",
    "1111100011011000",
    "1111000101110111",
    "1110101111011110",
    "1110100011100111",
    "1110100001111101",
    "1110100111000001",
    "1110101110111010",
    "1110110110111110",
    "1110111111000111",
    "1111001000110100",
    "1111010101000011",
    "1111100011100001",
    "1111110010000101",
    "1111111101011110",
    "1111111101000110",
    "1111111111001000",
    "1111110111110001",
    "1111101001111010",
    "1111011010100011",
    "1111001101000100",
    "1111000011110100",
    "1110111111111010",
    "1111000001100110",
    "1111001000110100",
    "1111010100110110",
    "1111100100101100",
    "1111110111001110",
    "1111110100011001",
    "1111011111001100",
    "1111001010010100",
    "1110110111101101",
    "1110101001001100",
    "1110100000001100",
    "1110011101010010",
    "1110100000100111",
    "1110101010000100",
    "1110111001010101",
    "1111001101101110",
    "1111100110001001",
    "1111111111010110",
    "1111100101011011",
    "1111001110111000",
    "1110111110001001",
    "1110110100100101",
    "1110110010010000",
    "1110110110001110",
    "1110111111001101",
    "1111001100001001",
    "1111011011111010",
    "1111101101000110",
    "1111111101111001",
    "1111110011110001",
    "1111101001111101",
    "1111100110000001",
    "1111101000010100",
    "1111101111110101",
    "1111111010011100",
    "1111111010001101",
    "1111110000000110",
    "1111101000001101",
    "1111100010101111",
    "1111011111011111",
    "1111011110010001",
    "1111011111101011",
    "1111100101101100",
    "1111110010110111",
    "1111110111011001",
    "1111011010010100",
    "1110111001101011",
    "1110011011000010",
    "1110000100000110",
    "1101111000110101",
    "1101111001111101",
    "1110000100111011",
    "1110010101001000",
    "1110100110000000",
    "1110110100011000",
    "1110111111001010",
    "1111000110101101",
    "1111001011111101",
    "1111010001010111",
    "1111011011000110",
    "1111101011110111",
    "1111111100101010",
    "1111100010001000",
    "1111001010100010",
    "1110111011011110",
    "1110111000110100",
    "1111000011100001",
    "1111011000000001",
    "1111110000001100",
    "1111111001010000",
    "1111100110100100",
    "1111010101110111",
    "1111000100010111",
    "1110110001000101",
    "1110011101110011",
    "1110001111011010",
    "1110001100001100",
    "1110011000011010",
    "1110110011111001",
    "1111011001010000",
    "1111111111101000",
    "1111100001110000",
    "1111010000011111",
    "1111001101000100",
    "1111010011111011",
    "1111011111101001",
    "1111101011001100",
    "1111110011001011",
    "1111110110101111",
    "1111110111010011",
    "1111110111010100",
    "1111111000110001",
    "1111111100011000",
    "1111111110101000",
    "1111111001010101",
    "1111110100001010",
    "1111101110101111",
    "1111101000001100",
    "1111011111101001",
    "1111010100110100",
    "1111001000011011",
    "1110111100001001",
    "1110110010000011",
    "1110101011101101",
    "1110101001111101",
    "1110101101001010",
    "1110110101010111",
    "1111000010011010",
    "1111010011000101",
    "1111100101001011",
    "1111110101101100",
    "1111111110011010",
    "1111111001011010",
    "1111111100000000",
    "1111111010100100",
    "1111101100010100",
    "1111011011010110",
    "1111001001011001",
    "1110110111010001",
    "1110100101100000",
    "1110010101010010",
    "1110001000100011",
    "1110000001101110",
    "1110000010010101",
    "1110001010100010",
    "1110011000101101",
    "1110101010010011",
    "1110111101010100",
    "1111010001110110",
    "1111101001100111",
    "1111111001111011",
    "1111011001011101",
    "1110111000101000",
    "1110011101000101",
    "1110001100100101",
    "1110001011000001",
    "1110011000110010",
    "1110110010110110",
    "1111010100100000",
    "1111111000100011",
    "1111100101010000",
    "1111000111111110",
    "1110110001100111",
    "1110100011011100",
    "1110011110001101",
    "1110100010101100",
    "1110110000111101",
    "1111000111110100",
    "1111100100100101",
    "1111111100110011",
    "1111100001001100",
    "1111001100100011",
    "1111000001010010",
    "1110111111111101",
    "1111000111110001",
    "1111010111001101",
    "1111101100100010",
    "1111111010010001",
    "1111011111110110",
    "1111000110111110",
    "1110110010010101",
    "1110100011110110",
    "1110011100011001",
    "1110011011111000",
    "1110100010000011",
    "1110101110111111",
    "1111000011001101",
    "1111011110101110",
    "1111111111101100",
    "1111011011000010",
    "1110110111100000",
    "1110011001101101",
    "1110000101011101",
    "1101111100010111",
    "1101111101011110",
    "1110000101110100",
    "1110010001111001",
    "1110011111000100",
    "1110101100100101",
    "1110111100100101",
    "1111010010011010",
    "1111101111111001",
    "1111101100100001",
    "1111001000010000",
    "1110101010001100",
    "1110011000011011",
    "1110010110001110",
    "1110100010011101",
    "1110111000000110",
    "1111010000101100",
    "1111100110110111",
    "1111111000000101",
    "1111111010110101",
    "1111101111100101",
    "1111100011111011",
    "1111010111010101",
    "1111001011111100",
    "1111000101100101",
    "1111001000001001",
    "1111010101101010",
    "1111101101000111",
    "1111110101100011",
    "1111011000001000",
    "1111000000000101",
    "1110110000111101",
    "1110101011110010",
    "1110101111011010",
    "1110111001011000",
    "1111000111010001",
    "1111011000111010",
    "1111110000000001",
    "1111110001111110",
    "1111001101111010",
    "1110100111100010",
    "1110000100111011",
    "1101101100001111",
    "1101100010000010",
    "1101100111100010",
    "1101111011001110",
    "1110011010000111",
    "1111000000011111",
    "1111101010010010",
    "1111101100110101",
    "1111001001100011",
    "1110101111110000",
    "1110100001101100",
    "1110011111010110",
    "1110100110001101",
    "1110110010001000",
    "1110111111000101",
    "1111001010000111",
    "1111010001111001",
    "1111010110100111",
    "1111011001011000",
    "1111011011100000",
    "1111011101110011",
    "1111100000101011",
    "1111100101001011",
    "1111101101100000",
    "1111111100001000",
    "1111101101110011",
    "1111010001111110",
    "1110110100101100",
    "1110011011100000",
    "1110001011000111",
    "1110000101101010",
    "1110001001110100",
    "1110010011110001",
    "1110011110111011",
    "1110100111110100",
    "1110101101101011",
    "1110110010010111",
    "1110111001001001",
    "1111000100101010",
    "1111010101011011",
    "1111101001001001",
    "1111111011101100",
    "1111110111010100",
    "1111110010101100",
    "1111110110010101",
    "1111111111110110",
    "1111110011111000",
    "1111100111010110",
    "1111011011101101",
    "1111010001100001",
    "1111001001011001",
    "1111000100011111",
    "1111000100010000",
    "1111001010000100",
    "1111010110100000",
    "1111101000101110",
    "1111111110001111",
    "1111101100100000",
    "1111011011010110",
    "1111010000111001",
    "1111001110000111",
    "1111010010001101",
    "1111011011100011",
    "1111101001101010",
    "1111111101100110",
    "1111100111100010",
    "1111000110100101",
    "1110100010111000",
    "1110000001101001",
    "1101101000010110",
    "1101011011000001",
    "1101011010101101",
    "1101100100111110",
    "1101110101000110",
    "1110000110010010",
    "1110010101000011",
    "1110100000110101",
    "1110101011111101",
    "1110111010011110",
    "1111001111011100",
    "1111101011010000",
    "1111110101001011",
    "1111010111001001",
    "1111000000000011",
    "1110110011111110",
    "1110110011111011",
    "1110111110000100",
    "1111001111000100",
    "1111100011010111",
    "1111110111110111",
    "1111110101111110",
    "1111101000100010",
    "1111100001011001",
    "1111100001001100",
    "1111100111101101",
    "1111110011110100",
    "1111111100100111",
    "1111101100010100",
    "1111011110000100",
    "1111010100010010",
    "1111010000100100",
    "1111010011010011",
    "1111011011110101",
    "1111101000101111",
    "1111111000001011",
    "1111110111111001",
    "1111101001101100",
    "1111011110110110",
    "1111011000010000",
    "1111010101100101",
    "1111010101011111",
    "1111010110000011",
    "1111010101100111",
    "1111010011100010",
    "1111010000011010",
    "1111001101111000",
    "1111001101110101",
    "1111010001111110",
    "1111011011001001",
    "1111101001001111",
    "1111111011001001",
    "1111110001010100",
    "1111011111000100",
    "1111010000111000",
    "1111001001000111",
    "1111001001011001",
    "1111010010101111",
    "1111100101001011",
    "1111111111000101",
    "1111100010100111",
    "1111000100001010",
    "1110101001111010",
    "1110010111100011",
    "1110001111000111",
    "1110010000010111",
    "1110011000111111",
    "1110100101100100",
    "1110110010100010",
    "1110111101011110",
    "1111000110001110",
    "1111001110101101",
    "1111011001011011",
    "1111100111111110",
    "1111111001111001",
    "1111110011000111",
    "1111100010010101",
    "1111010110100101",
    "1111010000111001",
    "1111001111111010",
    "1111010000100001",
    "1111001111100110",
    "1111001011000001",
    "1111000010011111",
    "1110110111100000",
    "1110101100011110",
    "1110100100000101",
    "1110100000010010",
    "1110100010001011",
    "1110101010001110",
    "1110111000001110",
    "1111001011001110",
    "1111100001001010",
    "1111110111000110",
    "1111110110010000",
    "1111101001101101",
    "1111100100101001",
    "1111100110011101",
    "1111101101001111",
    "1111110110111110",
    "1111111101000111",
    "1111101110110100",
    "1111011101100110",
    "1111001001111100",
    "1110110101110100",
    "1110100100010010",
    "1110011000100111",
    "1110010101000011",
    "1110011001110010",
    "1110100101010011",
    "1110110101111001",
    "1111001010100101",
    "1111100010110011",
    "1111111101101001",
    "1111100111000101",
    "1111001110111010",
    "1110111101111000",
    "1110110111011010",
    "1110111100101010",
    "1111001011110010",
    "1111100000111011",
    "1111110111111000",
    "1111110010011001",
    "1111011111011010",
    "1111001111100011",
    "1111000011001101",
    "1110111011011001",
    "1110111010000010",
    "1111000001001100",
    "1111010001100010",
    "1111101001111011",
    "1111111000110111",
    "1111011011011011",
    "1111000010010100",
    "1110110000110000",
    "1110100111111010",
    "1110100111001001",
    "1110101100110010",
    "1110110111000001",
    "1111000100010000",
    "1111010011010011",
    "1111100011010010",
    "1111110011001111",
    "1111111101110110",
    "1111110001001001",
    "1111100111011101",
    "1111100001000011",
    "1111011101110000",
    "1111011100111111",
    "1111011110001001",
    "1111100000110110",
    "1111100100111011",
    "1111101010001101",
    "1111110000001111",
    "1111110110000000",
    "1111111001111100",
    "1111111010011000",
    "1111110110001000",
    "1111101100111101",
    "1111011111110101",
    "1111010000011100",
    "1111000000111011",
    "1110110011001101",
    "1110101000111001",
    "1110100011001111",
    "1110100011000000",
    "1110101000001100",
    "1110110010000110",
    "1110111111010100",
    "1111001101111111",
    "1111011100001010",
    "1111101000011001",
    "1111110010001001",
    "1111111010000101",
    "1111111110010010",
    "1111110101101000",
    "1111101011010110",
    "1111100000000101",
    "1111010101011111",
    "1111001101101110",
    "1111001010101000",
    "1111001100111000",
    "1111010011110001",
    "1111011101011011",
    "1111100111101001",
    "1111110000111101",
    "1111111001100110",
    "1111111100110100",
    "1111110000101101",
    "1111100001100010",
    "1111010000110110",
    "1111000010000011",
    "1110111001010110",
    "1110111010010100",
    "1111000110011101",
    "1111011100000111",
    "1111110111000100",
    "1111101110000001",
    "1111011000000100",
    "1111001010000010",
    "1111000100110001",
    "1111000110111110",
    "1111001101110011",
    "1111010110010101",
    "1111011110011100",
    "1111100101110100",
    "1111101110001001",
    "1111111001111110",
    "1111110100110010",
    "1111011110001101",
    "1111000100011101",
    "1110101011001100",
    "1110010110100010",
    "1110001001100101",
    "1110000101010010",
    "1110001000000100",
    "1110001111000010",
    "1110010111000001",
    "1110011101110111",
    "1110100010101110",
    "1110100101101100",
    "1110100111100010",
    "1110101000111001",
    "1110101010000010",
    "1110101010101010",
    "1110101010101000",
    "1110101100101000",
    "1110110100111011",
    "1111000110000011",
    "1111011111100110",
    "1111111101001101",
    "1111100111100011",
    "1111010100101010",
    "1111001110001010",
    "1111010100011111",
    "1111100100011100",
    "1111111001100111",
    "1111110000001000",
    "1111011011111111",
    "1111001011101101",
    "1111000000110000",
    "1110111100011001",
    "1110111111010001",
    "1111001010000001",
    "1111011100100101",
    "1111110101100011",
    "1111101101101100",
    "1111010001000010",
    "1110111000110010",
    "1110101000011010",
    "1110100001011001",
    "1110100010111101",
    "1110101010110000",
    "1110110110000001",
    "1111000010001000",
    "1111001100111000",
    "1111010101111001",
    "1111011110110011",
    "1111101001111111",
    "1111111001010111",
    "1111110011000011",
    "1111011101111010",
    "1111001011001100",
    "1110111111000010",
    "1110111100010100",
    "1111000011010011",
    "1111010001111011",
    "1111100100110110",
    "1111111000100010",
    "1111110101110000",
    "1111101000000100",
    "1111011111101001",
    "1111011100101101",
    "1111011110101011",
    "1111100100100010",
    "1111101101000101",
    "1111110111001110",
    "1111111101111000",
    "1111110011010110",
    "1111101010000101",
    "1111100010110001",
    "1111011101101000",
    "1111011010011110",
    "1111011000111111",
    "1111011001001110",
    "1111011011010100",
    "1111011111010010",
    "1111100101000101",
    "1111101100100100",
    "1111110101101000",
    "1111111111111100",
    "1111110100011110",
    "1111101000001110",
    "1111011011101000",
    "1111001111010111",
    "1111000100100101",
    "1110111100101101",
    "1110111001010000",
    "1110111011100101",
    "1111000100010101",
    "1111010010111011",
    "1111100101011011",
    "1111111001000100",
    "1111110101010011",
    "1111101000100010",
    "1111100010011001",
    "1111100011101010",
    "1111101100011001",
    "1111111100001011",
    "1111101101101110",
    "1111010010111110",
    "1110110110000110",
    "1110011010100000",
    "1110000100001110",
    "1101110110110001",
    "1101110100000110",
    "1101111100000100",
    "1110001011111000",
    "1110011111101011",
    "1110110101000110",
    "1111001100100110",
    "1111100111101110",
    "1111111000110110",
    "1111010111000011",
    "1110110111001000",
    "1110011110011110",
    "1110010001110000",
    "1110010010101110",
    "1110011111000101",
    "1110110010111110",
    "1111001011100001",
    "1111100111001100",
    "1111111010100000",
    "1111011010101011",
    "1110111011110010",
    "1110100001000000",
    "1110001110001111",
    "1110000110011011",
    "1110001001101000",
    "1110010101010111",
    "1110100101110100",
    "1110110111110111",
    "1111001010001111",
    "1111011101010110",
    "1111110010000000",
    "1111110111100011",
    "1111100001001111",
    "1111001110011100",
    "1111000010011101",
    "1110111110111010",
    "1111000011000011",
    "1111001100000010",
    "1111010110010011",
    "1111011110111010",
    "1111100100101001",
    "1111100111111111",
    "1111101010110110",
    "1111101111110100",
    "1111111000111001",
    "1111111001101110",
    "1111101010001100",
    "1111011100011110",
    "1111010101010010",
    "1111011000010110",
    "1111100111010101",
    "1111111110111110",
    "1111011110010111",
    "1110111100000010",
    "1110011101100000",
    "1110000111011010",
    "1101111100101010",
    "1101111101110101",
    "1110001001001110",
    "1110011011011001",
    "1110110000011001",
    "1111000100110111",
    "1111010110101101",
    "1111100101110100",
    "1111110100010001",
    "1111111010110111",
    "1111100101101100",
    "1111001100100011",
    "1110110010011111",
    "1110011100000101",
    "1110001101101011",
    "1110001010000001",
    "1110010001010111",
    "1110100001111011",
    "1110111000111001",
    "1111010011010111",
    "1111101110110101",
    "1111110111000011",
    "1111100000111001",
    "1111010001000000",
    "1111001000111001",
    "1111001001001100",
    "1111010001100111",
    "1111100001000011",
    "1111110101101111",
    "1111110010100100",
    "1111011010111010",
    "1111000110011101",
    "1110111000001001",
    "1110110001111011",
    "1110110100011100",
    "1110111111001100",
    "1111010000011001",
    "1111100101001101",
    "1111111010011000",
    "1111110011000110",
    "1111100101011011",
    "1111011101101000",
    "1111011011100110",
    "1111011110100001",
    "1111100101001101",
    "1111101110101001",
    "1111111010001010",
    "1111111000011100",
    "1111101001010101",
    "1111011000101000",
    "1111000110101100",
    "1110110100010000",
    "1110100010100110",
    "1110010011010011",
    "1110001000000001",
    "1110000001110011",
    "1110000001000000",
    "1110000101010011",
    "1110001101111111",
    "1110011010010110",
    "1110101010110000",
    "1111000000000011",
    "1111011010100010",
    "1111111000111000",
    "1111101000000011",
    "1111001100110011",
    "1110111001111001",
    "1110110010011100",
    "1110110110101101",
    "1111000011111001",
    "1111010101001011",
    "1111100101011101",
    "1111110001001011",
    "1111110110110110",
    "1111111000001001",
    "1111111010001000",
    "1111111101011111",
    "1111101011111010",
    "1111010010011001",
    "1110110110001000",
    "1110011110000000",
    "1110010000000000",
    "1110001111011111",
    "1110011011110000",
    "1110110000110101",
    "1111001001101101",
    "1111100001101001",
    "1111110101001010",
    "1111111110000111",
    "1111111010000110",
    "1111111111110000",
    "1111110001001110",
    "1111011010011110",
    "1110111111011010",
    "1110100100111001",
    "1110001111110110",
    "1110000100001000",
    "1110000011011000",
    "1110001100011001",
    "1110011011101010",
    "1110101100101101",
    "1110111100000001",
    "1111001000110000",
    "1111010101010011",
    "1111100101010011",
    "1111111011001001",
    "1111101001011000",
    "1111001011101000",
    "1110110000011010",
    "1110011100010110",
    "1110010010001101",
    "1110010001011001",
    "1110010110011010",
    "1110011101000000",
    "1110100001111001",
    "1110100100000101",
    "1110100100110001",
    "1110100110001101",
    "1110101010010011",
    "1110110001110001",
    "1110111011110000",
    "1111000111011111",
    "1111010101001110",
    "1111100101101110",
    "1111111001001100",
    "1111110001100101",
    "1111011101101001",
    "1111001110101110",
    "1111000111110111",
    "1111001001110000",
    "1111010010001111",
    "1111011101001001",
    "1111100110100011",
    "1111101100001111",
    "1111101110101110",
    "1111110000101011",
    "1111110101010011",
    "1111111110110100",
    "1111110010101001",
    "1111100001011100",
    "1111010001000111",
    "1111000101001101",
    "1110111111111011",
    "1111000001011001",
    "1111000111111010",
    "1111010001000111",
    "1111011010111101",
    "1111100100011000",
    "1111101100111010",
    "1111110100001101",
    "1111111001101001",
    "1111111100011000",
    "1111111011110111",
    "1111111000001100",
    "1111110010101011",
    "1111101101011101",
    "1111101011000111",
    "1111101101101111",
    "1111110110010100",
    "1111111011110001",
    "1111101010101100",
    "1111011001010011",
    "1111001010010011",
    "1110111111010111",
    "1110111001000111",
    "1110110111010101",
    "1110111001010101",
    "1110111110010100",
    "1111000101011111",
    "1111001110010111",
    "1111011000110010",
    "1111100100111011",
    "1111110011010001",
    "1111111011110000",
    "1111101000010100",
    "1111010011010111",
    "1110111110101000",
    "1110101100000111",
    "1110011101110000",
    "1110010100110111",
    "1110010001111011",
    "1110010100101010",
    "1110011100100000",
    "1110101000111100",
    "1110111001101000",
    "1111001110000000",
    "1111100101000110",
    "1111111101001111",
    "1111101011100110",
    "1111010111100101",
    "1111001000100000",
    "1110111111011010",
    "1110111100011001",
    "1110111110101011",
    "1111000100110011",
    "1111001101000101",
    "1111010101101111",
    "1111011101000010",
    "1111100001110001",
    "1111100011011010",
    "1111100010100100",
    "1111100000110101",
    "1111100000001101",
    "1111100010010101",
    "1111100111101000",
    "1111101110111110",
    "1111110110001001",
    "1111111010100001",
    "1111111010011000",
    "1111110101101001",
    "1111101110001101",
    "1111100111011010",
    "1111100101000110",
    "1111101010011101",
    "1111111001011000",
    "1111101101111110",
    "1111001101101000",
    "1110101001001001",
    "1110000101010011",
    "1101100111001011",
    "1101010010111001",
    "1101001010110111",
    "1101001111001010",
    "1101011101011110",
    "1101110010100010",
    "1110001100010100",
    "1110101010001111",
    "1111001100001001",
    "1111110000110000",
    "1111101010111100",
    "1111001011100011",
    "1110110101101010",
    "1110101100111000",
    "1110110010000000",
    "1111000010111000",
    "1111011011101000",
    "1111110111111101",
    "1111101011100000",
    "1111010000111011",
    "1110111001011110",
    "1110100101101100",
    "1110010101101110",
    "1110001001100111",
    "1110000001000111",
    "1101111011011001",
    "1101110111100111",
    "1101110101000110",
    "1101110011100001",
    "1101110011000011",
    "1101110100001011",
    "1101110111100011",
    "1101111101000111",
    "1110000011110100",
    "1110001010001001",
    "1110001111000010",
    "1110010011100110",
    "1110011011001001",
    "1110101001010101",
    "1110111111110101",
    "1111011101001010",
    "1111111100111110",
    "1111100110001110",
    "1111010001001111",
    "1111000110001001",
    "1111000011011010",
    "1111000100111110",
    "1111000110010011",
    "1111000100011100",
    "1110111110110110",
    "1110110111011101",
    "1110110001110000",
    "1110110001100111",
    "1110111001010011",
    "1111001000000110",
    "1111011010101000",
    "1111101100000001",
    "1111110111101101",
    "1111111011000000",
    "1111110101101011",
    "1111101001111100",
    "1111011011010110",
    "1111001101110000",
    "1111000100010111",
    "1111000001001000",
    "1111000100111011",
    "1111010000010101",
    "1111100011100100",
    "1111111101110111",
    "1111100011000001",
    "1111000011001000",
    "1110100111011000",
    "1110010100010011",
    "1110001100110101",
    "1110010001000111",
    "1110011110010110",
    "1110110000000000",
    "1111000001011100",
    "1111001111100100",
    "1111011001011011",
    "1111011111101001",
    "1111100011101001",
    "1111100110110100",
    "1111101010001010",
    "1111101110101111",
    "1111110110011110",
    "1111111100010110",
    "1111101000110101",
    "1111010000000010",
    "1110110101101010",
    "1110011111000101",
    "1110010001101001",
    "1110010001000010",
    "1110011101011011",
    "1110110011010111",
    "1111001101100100",
    "1111100110110100",
    "1111111011100101",
    "1111110101010011",
    "1111101011100001",
    "1111100101100101",
    "1111100001110110",
    "1111011111011110",
    "1111011110000101",
    "1111011101011011",
    "1111011101001001",
    "1111011100100000",
    "1111011010101111",
    "1111010111101000",
    "1111010011110011",
    "1111010000100111",
    "1111001111101100",
    "1111010001111001",
    "1111010111001000",
    "1111011110010110",
    "1111100110000000",
    "1111101100101010",
    "1111110001101000",
    "1111110101000111",
    "1111111000001001",
    "1111111100011010",
    "1111111100010011",
    "1111110000101111",
    "1111100000100111",
    "1111001101000111",
    "1110111000101101",
    "1110100110101100",
    "1110011010010100",
    "1110010110001011",
    "1110011011101000",
    "1110101010100101",
    "1111000001010010",
    "1111011100110010",
    "1111111001010100",
    "1111101100110100",
    "1111011000110101",
    "1111001100111000",
    "1111001001111001",
    "1111001111101001",
    "1111011100111101",
    "1111110000001000",
    "1111111001000010",
    "1111100001001010",
    "1111001011000100",
    "1110111001010001",
    "1110101101101101",
    "1110101001001011",
    "1110101011010100",
    "1110110010101001",
    "1110111100111100",
    "1111000111101000",
    "1111010000011100",
    "1111010101011111",
    "1111010101101001",
    "1111010000101100",
    "1111000111010011",
    "1110111010110101",
    "1110101101001001",
    "1110100000010101",
    "1110010110101000",
    "1110010001111101",
    "1110010011101001",
    "1110011100000100",
    "1110101010001100",
    "1110111011110111",
    "1111001110000111",
    "1111011101110011",
    "1111101000011101",
    "1111101100101001",
    "1111101001111110",
    "1111100001001111",
    "1111010100011000",
    "1111000110000011",
    "1110111000111110",
    "1110101111100011",
    "1110101011001010",
    "1110101100001100",
    "1110110001100100",
    "1110111001111111",
    "1111000101000101",
    "1111010011101111",
    "1111100110111110",
    "1111111110100001",
    "1111100111110111",
    "1111010000000111",
    "1110111110011011",
    "1110110110001101",
    "1110111000011101",
    "1111000011000101",
    "1111010001111110",
    "1111100000100100",
    "1111101011101010",
    "1111110100001000",
    "1111111110110011",
    "1111101111010100",
    "1111010100010010",
    "1110110010110001",
    "1110010001100001",
    "1101111000001110",
    "1101101101000010",
    "1101110010000000",
    "1110000011011100",
    "1110011010101000",
    "1110110001000111",
    "1111000011010000",
    "1111010010000011",
    "1111100000110001",
    "1111110010000111",
    "1111111001011000",
    "1111100100110001",
    "1111010101011111",
    "1111010000110000",
    "1111011001100000",
    "1111101110100011",
    "1111110101011100",
    "1111011001011101",
    "1111000011010000",
    "1110110101110111",
    "1110110001011010",
    "1110110100110111",
    "1110111110110101",
    "1111001101111111",
    "1111100001001111",
    "1111110111011101",
    "1111110000111011",
    "1111011001111111",
    "1111000101111011",
    "1110110110101000",
    "1110101101001111",
    "1110101001101111",
    "1110101011110011",
    "1110110011001000",
    "1110111111101001",
    "1111010001000111",
    "1111100110101000",
    "1111111110010110",
    "1111101010011010",
    "1111010111000001",
    "1111001010000001",
    "1111000100101001",
    "1111000110100101",
    "1111001110110001",
    "1111011100001010",
    "1111101110001001",
    "1111111011101010",
    "1111100010001000",
    "1111000111000001",
    "1110101101000111",
    "1110010111100111",
    "1110001001011011",
    "1110000100010111",
    "1110001000011011",
    "1110010011101100",
    "1110100011010011",
    "1110110101001101",
    "1111001001010001",
    "1111100000010101",
    "1111111010110110",
    "1111101000101100",
    "1111001101111010",
    "1110111001010011",
    "1110101111000111",
    "1110110001010101",
    "1110111111000000",
    "1111010100101001",
    "1111101110000111",
    "1111111000000110",
    "1111100000000111",
    "1111001010110100",
    "1110111000110101",
    "1110101010111111",
    "1110100010100001",
    "1110100000111110",
    "1110100111110001",
    "1110110111100000",
    "1111001111010111",
    "1111101100011110",
    "1111110101011010",
    "1111011010111010",
    "1111000111101100",
    "1110111101110000",
    "1110111101001110",
    "1111000100100101",
    "1111010001010101",
    "1111100000100111",
    "1111110000001011",
    "1111111110101101",
    "1111110100001101",
    "1111101000100110",
    "1111011110010001",
    "1111010101000011",
    "1111001100101110",
    "1111000101000101",
    "1110111101110111",
    "1110110110110100",
    "1110110000000010",
    "1110101001111111",
    "1110100101101100",
    "1110100100001000",
    "1110100101110001",
    "1110101010010011",
    "1110110000101110",
    "1110110111111100",
    "1111000000001010",
    "1111001011111010",
    "1111011101110011",
    "1111110110100010",
    "1111101100000111",
    "1111001111010001",
    "1110111000101010",
    "1110101100111101",
    "1110101110000000",
    "1110111001011101",
    "1111001001111001",
    "1111011001101111",
    "1111100101111001",
    "1111101111010001",
    "1111111001010101",
    "1111111000100001",
    "1111100100111100",
    "1111001101101110",
    "1110110111100011",
    "1110100111110101",
    "1110100010101100",
    "1110101001010101",
    "1110111001111100",
    "1111010001001100",
    "1111101011011100",
    "1111111010000010",
    "1111100001011110",
    "1111001100111000",
    "1110111110011001",
    "1110110111101100",
    "1110111001101101",
    "1111000100001000",
    "1111010101010011",
    "1111101010101101",
    "1111111110110101",
    "1111101010101001",
    "1111011011010110",
    "1111010010110100",
    "1111010010010010",
    "1111011010000010",
    "1111101001011110",
    "1111111110100110",
    "1111101001101011",
    "1111010011000101",
    "1111000000110110",
    "1110110101011011",
    "1110110001100010",
    "1110110100011100",
    "1110111100110011",
    "1111001001101010",
    "1111011010101011",
    "1111101111110010",
    "1111110111101101",
    "1111011101101001",
    "1111000100011111",
    "1110101110111111",
    "1110011111000000",
    "1110010101011010",
    "1110010001111011",
    "1110010100000000",
    "1110011011000110",
    "1110100111000110",
    "1110110111111110",
    "1111001101010010",
    "1111100101101110",
    "1111111110100110",
    "1111101011100000",
    "1111011100000010",
    "1111010101010111",
    "1111011000100000",
    "1111100101001001",
    "1111111001100001",
    "1111101101000111",
    "1111010010000110",
    "1110111000101101",
    "1110100100000000",
    "1110010110010000",
    "1110010000110011",
    "1110010011011000",
    "1110011100011100",
    "1110101001100111",
    "1110111000010110",
    "1111000110101000",
    "1111010011001000",
    "1111011101011001",
    "1111100111000101",
    "1111110011010001",
    "1111111011011110",
    "1111100100111100",
    "1111001011111000",
    "1110110101010010",
    "1110100110010000",
    "1110100010100100",
    "1110101011010110",
    "1110111110100110",
    "1111011000110010",
    "1111110110000011",
    "1111101100110001",
    "1111010010001010",
    "1110111100010100",
    "1110101101011001",
    "1110100111010000",
    "1110101011000100",
    "1110111001010011",
    "1111010001001010",
    "1111110000100001",
    "1111101100001001",
    "1111001001100011",
    "1110101100001100",
    "1110010111011000",
    "1110001100011110",
    "1110001011000100",
    "1110010001010010",
    "1110011100011011",
    "1110101001011000",
    "1110110101011000",
    "1110111110101110",
    "1111000100101110",
    "1111000111111111",
    "1111001010000100",
    "1111001100111100",
    "1111010010010100",
    "1111011011011000",
    "1111101000100001",
    "1111111001010101",
    "1111110011011110",
    "1111100000000101",
    "1111001111000010",
    "1111000010111000",
    "1110111101001010",
    "1110111110001001",
    "1111000100110001",
    "1111001111111111",
    "1111011111001010",
    "1111110010001110",
    "1111110111001011",
    "1111011110100100",
    "1111000110110010",
    "1110110011010000",
    "1110100110111011",
    "1110100011010000",
    "1110100111111110",
    "1110110011000000",
    "1111000001101011",
    "1111010001100100",
    "1111100001101001",
    "1111110001111010",
    "1111111101000111",
    "1111101011010110",
    "1111011001101011",
    "1111001010000110",
    "1110111111001101",
    "1110111011100000",
    "1111000000001101",
    "1111001101001010",
    "1111100000110101",
    "1111111000110001",
    "1111101101101110",
    "1111010101100101",
    "1111000001011001",
    "1110110011010101",
    "1110101101000000",
    "1110101111001010",
    "1110111001110100",
    "1111001100001110",
    "1111100100101001",
    "1111111111101110",
    "1111100100101110",
    "1111001110000100",
    "1110111110110101",
    "1110111000101101",
    "1110111100000010",
    "1111000111101101",
    "1111011001111101",
    "1111110000101011",
    "1111110110100100",
    "1111011110100100",
    "1111001010001100",
    "1110111011111101",
    "1110110101010011",
    "1110110110100000",
    "1110111110101001",
    "1111001100001110",
    "1111011101100110",
    "1111110001011111",
    "1111111001010100",
    "1111100100001110",
    "1111010000110001",
    "1111000000100111",
    "1110110101010010",
    "1110101111111011",
    "1110110001000101",
    "1110111000010000",
    "1111000100010000",
    "1111010011011000",
    "1111100011110110",
    "1111110100000100",
    "1111111101000101",
    "1111110000100010",
    "1111100110111011",
    "1111100000110001",
    "1111011110100011",
    "1111100000100110",
    "1111100110111110",
    "1111110001010000",
    "1111111110010011",
    "1111110011101001",
    "1111100110111010",
    "1111011101100110",
    "1111011001010101",
    "1111011010011110",
    "1111100000000111",
    "1111101000010000",
    "1111110000010101",
    "1111110110001011",
    "1111111000011010",
    "1111110110110001",
    "1111110001111111",
    "1111101011010011",
    "1111100100000001",
    "1111011101000111",
    "1111010110111001",
    "1111010001000111",
    "1111001011001001",
    "1111000100101001",
    "1110111101101001",
    "1110110110100100",
    "1110110000001000",
    "1110101011000100",
    "1110100111110100",
    "1110100110100010",
    "1110100111001000",
    "1110101001011001",
    "1110101101010100",
    "1110110010110100",
    "1110111010001111",
    "1111000101010000",
    "1111010110110111",
    "1111110001001101",
    "1111101100001010",
    "1111000101000011",
    "1110011111011111",
    "1110000001111000",
    "1101110000111110",
    "1101101110011011",
    "1101110111100000",
    "1110000110110001",
    "1110010110010101",
    "1110100001111000",
    "1110101000000001",
    "1110101010010100",
    "1110101100000101",
    "1110110001000000",
    "1110111011001110",
    "1111001010101000",
    "1111011101010100",
    "1111110000110001",
    "1111111101000011",
    "1111101101000001",
    "1111011110110000",
    "1111010001100111",
    "1111000101011111",
    "1110111010111101",
    "1110110011000001",
    "1110101110100001",
    "1110101101111010",
    "1110110001000011",
    "1110110111000011",
    "1110111110100001",
    "1111000110010110",
    "1111001110100011",
    "1111011000010001",
    "1111100101000101",
    "1111110101100110",
    "1111110111000110",
    "1111100011101010",
    "1111010011010111",
    "1111001001001001",
    "1111000110011111",
    "1111001010101111",
    "1111010011101001",
    "1111011110011001",
    "1111101000011100",
    "1111101111111111",
    "1111110100000100",
    "1111110100101110",
    "1111110010100110",
    "1111101110101000",
    "1111101001100001",
    "1111100011110001",
    "1111011101011110",
    "1111010110011111",
    "1111001110101000",
    "1111000101111100",
    "1110111100110111",
    "1110110100001000",
    "1110101101001100",
    "1110101001100101",
    "1110101010011001",
    "1110101111101110",
    "1110111000101010",
    "1111000011101100",
    "1111001111001101",
    "1111011001101111",
    "1111100010001101",
    "1111100111111010",
    "1111101010010101",
    "1111101001000010",
    "1111100011111001",
    "1111011011000110",
    "1111001111011001",
    "1111000010000010",
    "1110110100100010",
    "1110101000010110",
    "1110011110101001",
    "1110010111111110",
    "1110010100010101",
    "1110010011011000",
    "1110010100100000",
    "1110010111011000",
    "1110011011111101",
    "1110100010011101",
    "1110101011000110",
    "1110110101111001",
    "1111000010101011",
    "1111010000111110",
    "1111100000011010",
    "1111110000010111",
    "1111111111101101",
    "1111110000011100",
    "1111100010010010",
    "1111010101101100",
    "1111001011000111",
    "1111000011001011",
    "1110111110001100",
    "1110111100010111",
    "1110111101101101",
    "1111000010000000",
    "1111001000111111",
    "1111010010010100",
    "1111011101001100",
    "1111101000101010",
    "1111110011011101",
    "1111111100010011",
    "1111111101110110",
    "1111111011101001",
    "1111111101010110",
    "1111111101001111",
    "1111110100111000",
    "1111101010110100",
    "1111100000110110",
    "1111011001010001",
    "1111010110100000",
    "1111011010110101",
    "1111100111110100",
    "1111111100110110",
    "1111101000110011",
    "1111001101101001",
    "1110110110100100",
    "1110100111011010",
    "1110100010000101",
    "1110100101110110",
    "1110101111110001",
    "1110111100001110",
    "1111001000001100",
    "1111010010111000",
    "1111011110001001",
    "1111101101010000",
    "1111111101010011",
    "1111100001101001",
    "1111000010111110",
    "1110100110110110",
    "1110010011000101",
    "1110001011111111",
    "1110010010101011",
    "1110100100100101",
    "1110111101001110",
    "1111010111011011",
    "1111101111001011",
    "1111111101111010",
    "1111110000111101",
    "1111101001110010",
    "1111100111100010",
    "1111101001001100",
    "1111101101101010",
    "1111110011100111",
    "1111111001110001",
    "1111111110111101",
    "1111111101011001",
    "1111111010110111",
    "1111110111110111",
    "1111110010001010",
    "1111100111111100",
    "1111011000101000",
    "1111000101010000",
    "1110110000010010",
    "1110011100110101",
    "1110001101110000",
    "1110000100110001",
    "1110000010010100",
    "1110000110010011",
    "1110010001001010",
    "1110100011010011",
    "1110111100001001",
    "1111011001001110",
    "1111110110000100",
    "1111110010011010",
    "1111100100110011",
    "1111100011010010",
    "1111101100101100",
    "1111111100110100",
    "1111110001100111",
    "1111100010111011",
    "1111011000101101",
    "1111010010001000",
    "1111001101001010",
    "1111001000010000",
    "1111000011001011",
    "1110111111100001",
    "1110111111100110",
    "1111000101101001",
    "1111010010101110",
    "1111100110001110",
    "1111111101111101",
    "1111101000111111",
    "1111010001011111",
    "1110111101100110",
    "1110101110111010",
    "1110100110011101",
    "1110100100100111",
    "1110101000101101",
    "1110110001011111",
    "1110111101001100",
    "1111001001110111",
    "1111010101101110",
    "1111011111011001",
    "1111100110010011",
    "1111101011010000",
    "1111110000011111",
    "1111111001000011",
    "1111111001000001",
    "1111100101110111",
    "1111010000000000",
    "1110111011100110",
    "1110101100101110",
    "1110100110000011",
    "1110100111100010",
    "1110101110011110",
    "1110110110111100",
    "1110111101011001",
    "1110111111111010",
    "1110111110011001",
    "1110111010001100",
    "1110110101000110",
    "1110110000111011",
    "1110101110100100",
    "1110101110000100",
    "1110101110110101",
    "1110110000000101",
    "1110110001011001",
    "1110110010101111",
    "1110110100100000",
    "1110110111001001",
    "1110111011010100",
    "1111000001110000",
    "1111001011000010",
    "1111010111001000",
    "1111100101000001",
    "1111110011000110",
    "1111111111001111",
    "1111111000010110",
    "1111110100110111",
    "1111110110010100",
    "1111111011111000",
    "1111111011101011",
    "1111110001100111",
    "1111100110011100",
    "1111011010010001",
    "1111001101000000",
    "1110111110101011",
    "1110101111111000",
    "1110100001111001",
    "1110010110110010",
    "1110010000100100",
    "1110010000011010",
    "1110010110001110",
    "1110100000111000",
    "1110101111110000",
    "1111000011101110",
    "1111011101110010",
    "1111111101101011",
    "1111011111000111",
    "1110111101010010",
    "1110100001111011",
    "1110010001001000",
    "1110001100011011",
    "1110010010000011",
    "1110011110101000",
    "1110101111001010",
    "1111000001111000",
    "1111010110010000",
    "1111101011101100",
    "1111111111100011",
    "1111101110011110",
    "1111100100101111",
    "1111100101111011",
    "1111110011011011",
    "1111110100010011",
    "1111010101100101",
    "1110110110010101",
    "1110011011111111",
    "1110001010001011",
    "1110000001110100",
    "1110000001101100",
    "1110000111110001",
    "1110010011001000",
    "1110100100011000",
    "1110111100011100",
    "1111011011001111",
    "1111111110100011",
    "1111011101111000",
    "1110111111000111",
    "1110101001010101",
    "1110011110100011",
    "1110011101110111",
    "1110100100011100",
    "1110101110101101",
    "1110111001110000",
    "1111000100010010",
    "1111001110000111",
    "1111010111110111",
    "1111100001111001",
    "1111101011111101",
    "1111110101001100",
    "1111111100111100",
    "1111111011010101",
    "1111101111111111",
    "1111011101110010",
    "1111000100010111",
    "1110100111001101",
    "1110001100101010",
    "1101111011000100",
    "1101110110011101",
    "1101111110111101",
    "1110010000001000",
    "1110100011010011",
    "1110110010111001",
    "1110111101010110",
    "1111000101110111",
    "1111010001100111",
    "1111100100001101",
    "1111111110000010",
    "1111100100100010",
    "1111001001101010",
    "1110110111001001",
    "1110110000000000",
    "1110110011001000",
    "1110111100000111",
    "1111000101101100",
    "1111001100010100",
    "1111001111101100",
    "1111010010010010",
    "1111010111110100",
    "1111100011010101",
    "1111110101011001",
    "1111110100010110",
    "1111011110011111",
    "1111001110000000",
    "1111000110101000",
    "1111001001011110",
    "1111010100101100",
    "1111100100011000",
    "1111110100010001",
    "1111111111011011",
    "1111111001011101",
    "1111111011010110",
    "1111111010100000",
    "1111101001011010",
    "1111010011101111",
    "1110111100101010",
    "1110100111010110",
    "1110010110010011",
    "1110001010110010",
    "1110000100110110",
    "1110000011100100",
    "1110000101110010",
    "1110001011000110",
    "1110010100001010",
    "1110100010100001",
    "1110110111011010",
    "1111010010101100",
    "1111110010011101",
    "1111101100111010",
    "1111001111110110",
    "1110111001110111",
    "1110101100100101",
    "1110100111101101",
    "1110101001111100",
    "1110110010001000",
    "1110111111110101",
    "1111010011001000",
    "1111101011110100",
    "1111110111001111",
    "1111011000101000",
    "1110111011111010",
    "1110100100110100",
    "1110010110001001",
    "1110010000110110",
    "1110010100000000",
    "1110011101010111",
    "1110101010100010",
    "1110111001101011",
    "1111001001111100",
    "1111011010111100",
    "1111101100010001",
    "1111111100111010",
    "1111110100111100",
    "1111101011011110",
    "1111101000010100",
    "1111101100001010",
    "1111110110101111",
    "1111111001001001",
    "1111100101101010",
    "1111010001101001",
    "1111000000000010",
    "1110110011101100",
    "1110101110101110",
    "1110110010100010",
    "1110111111110110",
    "1111010110010010",
    "1111110100010000",
    "1111101001001111",
    "1111000110011000",
    "1110100111101000",
    "1110010000111011",
    "1110000100101110",
    "1110000011100001",
    "1110001011101010",
    "1110011010111000",
    "1110110000011100",
    "1111001100111111",
    "1111110000100011",
    "1111100110101001",
    "1110111101000000",
    "1110011000001001",
    "1101111101010001",
    "1101110000000011",
    "1101110000110000",
    "1101111011111111",
    "1110001100110000",
    "1110011110010001",
    "1110101101100000",
    "1110111001110101",
    "1111000100000001",
    "1111001101011011",
    "1111010111000011",
    "1111100000111110",
    "1111101010101110",
    "1111110011111010",
    "1111111100101011",
    "1111111010000011",
    "1111101111000011",
    "1111100001100100",
    "1111010010010010",
    "1111000011000101",
    "1110110110000011",
    "1110101100100011",
    "1110100110110100",
    "1110100100001011",
    "1110100011011101",
    "1110100011100100",
    "1110100011111000",
    "1110100100101001",
    "1110100110110111",
    "1110101011110111",
    "1110110100011101",
    "1111000000110000",
    "1111001111111000",
    "1111100000010101",
    "1111110000011010",
    "1111111110100100",
    "1111110110000110",
    "1111101101111001",
    "1111101000101000",
    "1111100101111011",
    "1111100101000110",
    "1111100101010101",
    "1111100101101001",
    "1111100101001110",
    "1111100011110110",
    "1111100001101011",
    "1111011111001000",
    "1111011100100001",
    "1111011001111010",
    "1111010111000110",
    "1111010011111100",
    "1111010000101100",
    "1111001101111011",
    "1111001100110010",
    "1111001110100100",
    "1111010100011100",
    "1111011110101001",
    "1111101100100011",
    "1111111100101010",
    "1111110010111100",
    "1111100100001011",
    "1111011000101100",
    "1111010001100001",
    "1111001111000111",
    "1111010001010111",
    "1111010111101111",
    "1111100001011010",
    "1111101101001101",
    "1111111001110011",
    "1111111010000110",
    "1111101111111010",
    "1111101000101111",
    "1111100101101010",
    "1111100111101001",
    "1111101111000110",
    "1111111011110001",
    "1111110011010001",
    "1111011111101000",
    "1111001011000111",
    "1110110111100011",
    "1110100110011011",
    "1110011000011110",
    "1110001110000111",
    "1110000111011101",
    "1110000100110001",
    "1110000110011111",
    "1110001101000000",
    "1110011000011110",
    "1110101000010011",
    "1110111010101111",
    "1111001101000000",
    "1111011011110111",
    "1111100100010101",
    "1111100100110011",
    "1111011101011001",
    "1111010000001010",
    "1111000000010101",
    "1110110001101001",
    "1110100111010101",
    "1110100011101001",
    "1110100111011101",
    "1110110010010111",
    "1111000011001010",
    "1111011000000100",
    "1111101111010101",
    "1111111000101101",
    "1111100001011100",
    "1111001011110101",
    "1110111000011101",
    "1110100111100010",
    "1110011001001100",
    "1110001101101000",
    "1110000101011010",
    "1110000001000111",
    "1110000001010000",
    "1110000101111100",
    "1110001110101000",
    "1110011010001100",
    "1110100111000110",
    "1110110100001011",
    "1111000001111101",
    "1111010010011010",
    "1111100111100001",
    "1111111110011111",
    "1111100010000000",
    "1111000111101111",
    "1110110101010111",
    "1110101111110110",
    "1110111001010101",
    "1111001111101100",
    "1111101101011000",
    "1111110100110010",
    "1111011101010100",
    "1111010000001100",
    "1111001110101011",
    "1111010111100101",
    "1111101000001000",
    "1111111101000101",
    "1111101100101010",
    "1111011000001000",
    "1111001000000100",
    "1110111111000111",
    "1110111111011100",
    "1111001010001011",
    "1111011110001101",
    "1111111000010001",
    "1111101100100001",
    "1111010101001000",
    "1111000101000001",
    "1110111101111010",
    "1110111111101001",
    "1111001000100111",
    "1111010110101000",
    "1111100111110111",
    "1111111010100100",
    "1111110010111100",
    "1111100010110100",
    "1111010111100111",
    "1111010011101010",
    "1111011000010001",
    "1111100100110110",
    "1111110110110011",
    "1111110101100001",
    "1111100011111011",
    "1111010111000011",
    "1111001111110011",
    "1111001101011100",
    "1111001110001001",
    "1111010000000010",
    "1111010010000010",
    "1111010100101100",
    "1111011010010011",
    "1111100101110001",
    "1111111001000101",
    "1111101100001111",
    "1111001101100001",
    "1110101111110001",
    "1110011000010000",
    "1110001010110100",
    "1110001000100000",
    "1110001111101001",
    "1110011100110010",
    "1110101011111111",
    "1110111010001111",
    "1111000110010010",
    "1111010000110101",
    "1111011011110101",
    "1111101000100111",
    "1111110110101000",
    "1111111100101101",
    "1111110101001110",
    "1111110110010110",
    "1111111110001001",
    "1111101001100001",
    "1111001111101011",
    "1110110101101110",
    "1110100000011001",
    "1110010010111101",
    "1110001110010110",
    "1110010001100110",
    "1110011010001111",
    "1110100101011101",
    "1110110000111001",
    "1110111011010001",
    "1111000100100000",
    "1111001101001110",
    "1111010110000110",
    "1111011111011110",
    "1111101001000010",
    "1111110010000110",
    "1111111001110010",
    "1111111111001001",
    "1111111110010110",
    "1111111110110001",
    "1111111110110010",
    "1111111011111101",
    "1111111010011111",
    "1111111011101001",
    "1111111111111011",
    "1111111000111011",
    "1111101111100101",
    "1111100100101110",
    "1111011000111001",
    "1111001100101010",
    "1111000000110000",
    "1110110110010000",
    "1110101110011110",
    "1110101010110000",
    "1110101100001110",
    "1110110011000110",
    "1110111110101110",
    "1111001101001111",
    "1111011100000101",
    "1111101000110000",
    "1111110001011110",
    "1111110101101100",
    "1111110110000010",
    "1111110011111111",
    "1111110001010000",
    "1111101111001001",
    "1111101110000111",
    "1111101101110101",
    "1111101101011100",
    "1111101011111010",
    "1111101000100010",
    "1111100011001111",
    "1111011100101000",
    "1111010101110010",
    "1111010000000011",
    "1111001100101101",
    "1111001100110011",
    "1111010001001100",
    "1111011010001111",
    "1111100111110100",
    "1111111000110101",
    "1111110100100001",
    "1111100010110110",
    "1111010100101001",
    "1111001100000010",
    "1111001010011001",
    "1111010000000111",
    "1111011100110111",
    "1111101111101110",
    "1111111000111011",
    "1111011111101011",
    "1111000111011111",
    "1110110011010101",
    "1110100101011000",
    "1110011110100110",
    "1110011110101110",
    "1110100100100010",
    "1110101110011001",
    "1110111010110111",
    "1111001000110100",
    "1111010111001001",
    "1111100100011101",
    "1111101111000011",
    "1111110101010001",
    "1111110110010111",
    "1111110010111000",
    "1111101100111111",
    "1111101000001010",
    "1111101000001001",
    "1111101111100101",
    "1111111110110010",
    "1111101100011011",
    "1111010110001000",
    "1111000010100111",
    "1110110101001000",
    "1110101110111011",
    "1110101111010001",
    "1110110100100111",
    "1110111110000101",
    "1111001011110111",
    "1111011110001101",
    "1111110100100100",
    "1111110011010000",
    "1111011100101110",
    "1111001011011000",
    "1111000001101100",
    "1111000000001111",
    "1111000101101010",
    "1111001111111111",
    "1111011101110111",
    "1111101111000100",
    "1111111100000010",
    "1111100100000000",
    "1111001010110100",
    "1110110011110110",
    "1110100011000101",
    "1110011011011000",
    "1110011101011100",
    "1110100111100101",
    "1110110110010011",
    "1111000110001110",
    "1111010101101010",
    "1111100101001001",
    "1111110110011010",
    "1111110101011100",
    "1111011111100011",
    "1111001011011001",
    "1110111101111010",
    "1110111011100001",
    "1111000110010000",
    "1111011100101110",
    "1111111010100111",
    "1111100101110100",
    "1111001001111101",
    "1110110101010000",
    "1110101000111110",
    "1110100100011111",
    "1110100110001000",
    "1110101011110101",
    "1110110011110001",
    "1110111100100101",
    "1111000101100111",
    "1111001111001100",
    "1111011010011101",
    "1111101000100101",
    "1111111010000110",
    "1111110001101110",
    "1111011101001001",
    "1111001011001100",
    "1110111110111111",
    "1110111010011101",
    "1110111101100110",
    "1111000110100101",
    "1111010010100001",
    "1111011110011111",
    "1111101000011010",
    "1111101111001110",
    "1111110010111010",
    "1111110011111110",
    "1111110010110110",
    "1111101111100010",
    "1111101001101101",
    "1111100001010000",
    "1111010110101100",
    "1111001011011001",
    "1111000001100110",
    "1110111011100101",
    "1110111011010100",
    "1111000001110000",
    "1111001110101000",
    "1111100000011111",
    "1111110100111111",
    "1111110110101110",
    "1111100101010011",
    "1111011000100011",
    "1111010001000111",
    "1111001110011100",
    "1111001111010001",
    "1111010001111101",
    "1111010101001101",
    "1111011000010001",
    "1111011011000100",
    "1111011110000100",
    "1111100010010100",
    "1111101001010110",
    "1111110100110100",
    "1111111010011100",
    "1111100101001101",
    "1111001101111000",
    "1110110111111110",
    "1110100110111110",
    "1110011101011001",
    "1110011011111100",
    "1110100001011111",
    "1110101100000010",
    "1110111001011011",
    "1111001000000001",
    "1111010110101101",
    "1111100100100010",
    "1111110000000110",
    "1111110111011011",
    "1111111000010001",
    "1111110001000000",
    "1111100001100110",
    "1111001100000010",
    "1110110011111011",
    "1110011101101110",
    "1110001101010110",
    "1110000101001000",
    "1110000101001011",
    "1110001011100101",
    "1110010101011011",
    "1110011111111101",
    "1110101001000100",
    "1110110000001000",
    "1110110110000100",
    "1110111100110101",
    "1111000110101010",
    "1111010100111011",
    "1111100111101101",
    "1111111101110011",
    "1111101011000010",
    "1111010101101100",
    "1111000100100010",
    "1110111001000100",
    "1110110011110100",
    "1110110100010011",
    "1110111001010001",
    "1111000000111101",
    "1111001001011001",
    "1111010001000101",
    "1111010111001101",
    "1111011101000101",
    "1111100101111100",
    "1111110100101000",
    "1111110101111111",
    "1111011100011001",
    "1111000011101111",
    "1110110001110110",
    "1110101011010011",
    "1110110001110001",
    "1111000010111011",
    "1111011001111101",
    "1111110001101010",
    "1111111001100111",
    "1111101001000101",
    "1111011100001110",
    "1111010010001101",
    "1111001010110100",
    "1111000110111111",
    "1111001000011101",
    "1111010000011111",
    "1111011111000111",
    "1111110010101010",
    "1111111000000000",
    "1111100100010011",
    "1111010100101100",
    "1111001010001100",
    "1111000100101001",
    "1111000011101001",
    "1111000110110111",
    "1111001110010010",
    "1111011001110010",
    "1111101000110001",
    "1111111001111110",
    "1111110100100010",
    "1111100101011000",
    "1111011011010011",
    "1111011000011011",
    "1111011101101001",
    "1111101010010101",
    "1111111100010101",
    "1111101111010001",
    "1111011011110000",
    "1111001011101010",
    "1111000000011111",
    "1110111010100011",
    "1110111001011011",
    "1110111100010011",
    "1111000011000001",
    "1111001110101011",
    "1111100000111110",
    "1111111010111011",
    "1111100100001110",
    "1110111111110011",
    "1110011100100110",
    "1101111111111011",
    "1101101101110011",
    "1101100111010000",
    "1101101010010011",
    "1101110011000000",
    "1101111101001100",
    "1110000101111110",
    "1110001100100110",
    "1110010011011000",
    "1110011110101110",
    "1110110010010000",
    "1111001110101011",
    "1111110000110011",
    "1111101101011100",
    "1111010010110001",
    "1111000100010010",
    "1111000011101010",
    "1111001110010110",
    "1111011111010111",
    "1111110001010011",
    "1111111111111011",
    "1111110110101010",
    "1111110010011011",
    "1111110001111010",
    "1111110011001001",
    "1111110100101101",
    "1111110110010010",
    "1111111000001100",
    "1111111011001111",
    "1111111111111011",
    "1111111001011110",
    "1111110010000110",
    "1111101010110011",
    "1111100100100111",
    "1111100000011001",
    "1111011110111010",
    "1111100000011110",
    "1111100100110110",
    "1111101011100010",
    "1111110100010001",
    "1111111111011111",
    "1111110001101111",
    "1111011110100100",
    "1111000111010101",
    "1110101110001111",
    "1110010110111110",
    "1110000101110100",
    "1101111110011011",
    "1110000011001010",
    "1110010100101111",
    "1110110010000000",
    "1111010111100000",
    "1111111111111100",
    "1111011010110000",
    "1110111101111101",
    "1110101100101101",
    "1110100111100000",
    "1110101100000101",
    "1110110110100111",
    "1111000010111101",
    "1111001110000111",
    "1111010110101111",
    "1111011101001110",
    "1111100011011101",
    "1111101011101111",
    "1111110111101010",
    "1111111000101111",
    "1111100111001101",
    "1111010110000011",
    "1111000111011010",
    "1110111100010111",
    "1110110100100111",
    "1110101111000010",
    "1110101010011101",
    "1110100110100000",
    "1110100011101111",
    "1110100011001111",
    "1110100110001001",
    "1110101101010010",
    "1110111000101101",
    "1111000111011011",
    "1111010111110101",
    "1111101000001011",
    "1111110110110111",
    "1111111101001000",
    "1111110100010101",
    "1111101110110101",
    "1111101100100111",
    "1111101101010101",
    "1111110000011001",
    "1111110100111001",
    "1111111010000101",
    "1111111111101000",
    "1111111010001111",
    "1111110011001010",
    "1111101010110111",
    "1111100001101001",
    "1111011000010101",
    "1111001111111011",
    "1111001001001110",
    "1111000100011100",
    "1111000001010100",
    "1110111111000111",
    "1110111100111010",
    "1110111001111010",
    "1110110101011101",
    "1110101111010010",
    "1110100111100010",
    "1110011110101000",
    "1110010101001110",
    "1110001100010110",
    "1110000101001000",
    "1110000000110000",
    "1110000000001101",
    "1110000100000110",
    "1110001100101101",
    "1110011010001111",
    "1110101100111000",
    "1111000100011111",
    "1111100000000101",
    "1111111101110000",
    "1111100101010011",
    "1111001100001001",
    "1110111000110010",
    "1110101011110111",
    "1110100100010101",
    "1110100000001100",
    "1110011101010110",
    "1110011010011000",
    "1110010110111011",
    "1110010011100010",
    "1110010001001111",
    "1110010000110101",
    "1110010010101001",
    "1110010110011111",
    "1110011011110111",
    "1110100010010000",
    "1110101001011101",
    "1110110001011010",
    "1110111010010110",
    "1111000100010111",
    "1111001111011110",
    "1111011011101011",
    "1111101001001001",
    "1111111000001001",
    "1111110111000011",
    "1111100100110001",
    "1111010001111000",
    "1110111111111011",
    "1110110000101011",
    "1110100101100111",
    "1110011111011100",
    "1110011110000010",
    "1110100000011010",
    "1110100101010010",
    "1110101011011001",
    "1110110010000011",
    "1110111001000110",
    "1111000000110110",
    "1111001001100101",
    "1111010011010000",
    "1111011101100000",
    "1111100111110001",
    "1111110010001010",
    "1111111101111001",
    "1111110011010010",
    "1111100000011010",
    "1111001001111101",
    "1110110010011010",
    "1110011101100011",
    "1110001111001101",
    "1110001001111111",
    "1110001110011011",
    "1110011011010001",
    "1110101110100100",
    "1111000110011010",
    "1111100001001101",
    "1111111101010100",
    "1111100111010001",
    "1111001111001010",
    "1110111100111000",
    "1110110010011100",
    "1110110000101110",
    "1110110111010000",
    "1111000100101111",
    "1111010111100010",
    "1111101110000000",
    "1111111001100011",
    "1111100001001010",
    "1111001010111101",
    "1110111001011000",
    "1110101110101001",
    "1110101100010011",
    "1110110010110011",
    "1111000001000101",
    "1111010100100010",
    "1111101001101100",
    "1111111101000001",
    "1111110100001101",
    "1111101011100110",
    "1111101001001011",
    "1111101011111101",
    "1111110010010100",
    "1111111010100011",
    "1111111100101101",
    "1111110100101100",
    "1111101110010001",
    "1111101010000111",
    "1111101000101100",
    "1111101001110011",
    "1111101100110001",
    "1111110000010101",
    "1111110011000100",
    "1111110011110001",
    "1111110001110111",
    "1111101101101100",
    "1111101000011101",
    "1111100011110110",
    "1111100001011111",
    "1111100010011101",
    "1111100111001010",
    "1111101111010101",
    "1111111010010100",
    "1111111000110111",
    "1111101011101001",
    "1111011111110000",
    "1111010110111111",
    "1111010010111011",
    "1111010100011010",
    "1111011011010100",
    "1111100110100101",
    "1111110100011001",
    "1111111101001100",
    "1111101111110110",
    "1111100100001110",
    "1111011001101011",
    "1111001110100110",
    "1111000000111101",
    "1110101111101100",
    "1110011011101000",
    "1110000111010001",
    "1101110101111100",
    "1101101010101011",
    "1101100110111100",
    "1101101010010110",
    "1101110010111001",
    "1101111110000010",
    "1110001001110100",
    "1110010101101100",
    "1110100010010101",
    "1110110000111001",
    "1111000010000011",
    "1111010101010010",
    "1111101000111001",
    "1111111010110001",
    "1111110110111100",
    "1111101101001110",
    "1111100111101111",
    "1111100101010111",
    "1111100100110001",
    "1111100101000101",
    "1111100110001101",
    "1111101000010101",
    "1111101011101111",
    "1111110000011001",
    "1111110101111111",
    "1111111011111000",
    "1111111110101000",
    "1111111010011001",
    "1111110111110110",
    "1111110111000011",
    "1111110111100001",
    "1111111000011000",
    "1111111000100010",
    "1111110110111000",
    "1111110010101000",
    "1111101011100101",
    "1111100010010100",
    "1111011000000011",
    "1111001110010111",
    "1111000110101111",
    "1111000010001101",
    "1111000001010100",
    "1111000100000110",
    "1111001010011101",
    "1111010011111100",
    "1111100000001101",
    "1111101110101001",
    "1111111110011010",
    "1111110001100110",
    "1111100010101001",
    "1111010101101100",
    "1111001011011000",
    "1111000011111000",
    "1110111110111101",
    "1110111100001110",
    "1110111011010100",
    "1110111100001001",
    "1110111110111101",
    "1111000100100101",
    "1111001110011110",
    "1111011110000101",
    "1111110011110000",
    "1111110001110010",
    "1111010101111011",
    "1110111100111100",
    "1110101010111100",
    "1110100010011101",
    "1110100011100010",
    "1110101011110011",
    "1110110111101000",
    "1111000011011010",
    "1111001100110010",
    "1111010010110001",
    "1111010101010111",
    "1111010100110001",
    "1111010001000101",
    "1111001010000111",
    "1111000000001000",
    "1110110100001101",
    "1110101000011110",
    "1110011111101011",
    "1110011100000101",
    "1110011110110101",
    "1110100111001011",
    "1110110011000001",
    "1110111111101000",
    "1111001010110010",
    "1111010011100111",
    "1111011011010100",
    "1111100100110100",
    "1111110010111001",
    "1111111001001110",
    "1111100000111001",
    "1111000111100000",
    "1110110001010100",
    "1110100010000010",
    "1110011011011000",
    "1110011100001111",
    "1110100001100110",
    "1110101000000100",
    "1110101101010110",
    "1110110000110000",
    "1110110010111101",
    "1110110101000011",
    "1110110111110111",
    "1110111011011110",
    "1110111111010100",
    "1111000011101001",
    "1111001010011011",
    "1111010110000110",
    "1111100111111110",
    "1111111110110010",
    "1111101001011001",
    "1111010101110111",
    "1111001011010001",
    "1111001011101111",
    "1111010101110110",
    "1111100101110100",
    "1111110111110100",
    "1111110110001111",
    "1111100100000110",
    "1111010000010111",
    "1110111010011011",
    "1110100011010101",
    "1110001101111011",
    "1101111110000100",
    "1101110110101000",
    "1101111000110000",
    "1110000011100100",
    "1110010101010010",
    "1110101100010100",
    "1111000111011000",
    "1111100101001011",
    "1111111100010111",
    "1111100000011100",
    "1111001010100000",
    "1110111101001111",
    "1110111001001011",
    "1110111100010001",
    "1111000011000001",
    "1111001010000001",
    "1111001111011010",
    "1111010011011000",
    "1111010111011111",
    "1111011101010100",
    "1111100101010011",
    "1111101110001110",
    "1111110101011110",
    "1111111000011101",
    "1111110101101100",
    "1111101101101100",
    "1111100010110011",
    "1111011000011010",
    "1111010001100110",
    "1111010000010100",
    "1111010101001110",
    "1111100000000010",
    "1111110000010001",
    "1111111010101101",
    "1111100001111110",
    "1111000111000001",
    "1110101011111100",
    "1110010010111110",
    "1101111110001101",
    "1101101111000000",
    "1101100101110001",
    "1101100001111101",
    "1101100010101100",
    "1101100111101101",
    "1101110010010010",
    "1110000100011000",
    "1110011111001101",
    "1111000001111000",
    "1111101000101001",
    "1111110001111111",
    "1111010011101100",
    "1111000000010100",
    "1110111000101000",
    "1110111010010011",
    "1111000001011100",
    "1111001010010001",
    "1111010010100010",
    "1111011001110100",
    "1111100000110011",
    "1111101000100010",
    "1111110001100010",
    "1111111011010111",
    "1111111011010110",
    "1111110100101111",
    "1111110010110001",
    "1111110110101111",
    "1111111111001110",
    "1111110000010000",
    "1111011110010111",
    "1111001100100001",
    "1110111110000100",
    "1110110101111100",
    "1110110101110010",
    "1110111101011011",
    "1111001010110100",
    "1111011011000010",
    "1111101100011100",
    "1111111111111001",
    "1111100111111111",
    "1111001010110101",
    "1110101010001111",
    "1110001010111100",
    "1101110010110110",
    "1101100111010001",
    "1101101010101101",
    "1101111011000111",
    "1110010010110110",
    "1110101011010110",
    "1110111111000111",
    "1111001100000111",
    "1111010101000110",
    "1111011111001111",
    "1111101111001000",
    "1111111001111100",
    "1111011111100110",
    "1111001000010011",
    "1110111010110101",
    "1110111011100101",
    "1111001010100000",
    "1111100011000011",
    "1111111111001000",
    "1111100110011111",
    "1111010000110011",
    "1111000000001000",
    "1110110011101001",
    "1110101001101000",
    "1110100000100011",
    "1110010111111110",
    "1110010000011010",
    "1110001010111010",
    "1110001000100010",
    "1110001001101111",
    "1110001110000000",
    "1110010100100100",
    "1110011100011100",
    "1110100101111001",
    "1110110010011010",
    "1111000011101111",
    "1111011010110100",
    "1111110110011110",
    "1111101100100100",
    "1111010010110011",
    "1111000000011001",
    "1110110111111100",
    "1110111001010011",
    "1111000001101100",
    "1111001101010001",
    "1111011000101010",
    "1111100010010100",
    "1111101010011110",
    "1111110010011001",
    "1111111011001111",
    "1111111010111100",
    "1111110001100110",
    "1111101010101010",
    "1111100111111011",
    "1111101010100110",
    "1111110010111011",
    "1111111111111000",
    "1111101111101100",
    "1111011111000000",
    "1111010000011001",
    "1111000110010110",
    "1111000010111001",
    "1111000111010000",
    "1111010011011100",
    "1111100110000110",
    "1111111100100111",
    "1111101100001100",
    "1111010111011010",
    "1111000111001001",
    "1110111100100001",
    "1110111000000001",
    "1110111001111101",
    "1111000011000110",
    "1111010100011000",
    "1111101110000110",
    "1111110001010000",
    "1111001101011100",
    "1110101011100110",
    "1110010000110001",
    "1110000000010001",
    "1101111010101011",
    "1101111101111010",
    "1110000110001110",
    "1110010000000101",
    "1110011001101010",
    "1110100011010011",
    "1110101111000101",
    "1110111110111011",
    "1111010011010111",
    "1111101010101110",
    "1111111110011001",
    "1111101100000100",
    "1111100001011100",
    "1111011111111111",
    "1111100111000101",
    "1111110100100100",
    "1111111010010011",
    "1111101000010101",
    "1111010111110001",
    "1111001010010011",
    "1111000001001000",
    "1110111100111111",
    "1110111110011100",
    "1111000110000001",
    "1111010011111011",
    "1111100111101101",
    "1111111111111100",
    "1111100110000001",
    "1111001101101000",
    "1110111010000001",
    "1110101101010001",
    "1110101000000110",
    "1110101001110111",
    "1110110000111101",
    "1110111011010100",
    "1111000111001011",
    "1111010100000000",
    "1111100010110110",
    "1111110101100111",
    "1111110010011111",
    "1111010110011000",
    "1110111001001100",
    "1110011111011110",
    "1110001101110011",
    "1110000111000100",
    "1110001011100011",
    "1110011000111010",
    "1110101011101011",
    "1111000001000010",
    "1111010111111100",
    "1111110000100101",
    "1111110101000100",
    "1111011010011101",
    "1111000010110110",
    "1110110010110110",
    "1110101111001010",
    "1110111010111000",
    "1111010101101001",
    "1111111011010001",
    "1111011010111101",
    "1110110100011101",
    "1110010110111011",
    "1110000101010010",
    "1101111111101110",
    "1110000100100100",
    "1110010001101110",
    "1110100110000000",
    "1111000000100011",
    "1111100000001000",
    "1111111101110001",
    "1111011101000111",
    "1111000001111110",
    "1110101111011001",
    "1110100110001101",
    "1110100100110100",
    "1110100111111100",
    "1110101100000111",
    "1110101110111010",
    "1110101111100001",
    "1110101110100011",
    "1110101101010010",
    "1110101100111000",
    "1110101101101101",
    "1110101111100011",
    "1110110001110001",
    "1110110011110100",
    "1110110101010011",
    "1110110101111100",
    "1110110110000011",
    "1110110110111110",
    "1110111010111101",
    "1111000100000101",
    "1111010011010000",
    "1111100111110011",
    "1111111111001101",
    "1111101010001100",
    "1111011000011101",
    "1111001110010001",
    "1111001100000111",
    "1111010000100100",
    "1111011001001110",
    "1111100011100001",
    "1111101101011001",
    "1111110101100100",
    "1111111011011001",
    "1111111110101101",
    "1111111111100111",
    "1111111110000101",
    "1111111001110110",
    "1111110010100011",
    "1111100111111111",
    "1111011010101010",
    "1111001100000001",
    "1110111110010010",
    "1110110011111110",
    "1110101111011100",
    "1110110010011010",
    "1110111101011100",
    "1111001111011100",
    "1111100101110110",
    "1111111101010011",
    "1111101101011100",
    "1111011101000101",
    "1111010011000001",
    "1111001111100110",
    "1111010010011111",
    "1111011011010001",
    "1111101001101000",
    "1111111101000011",
    "1111101011110110",
    "1111010011100110",
    "1110111101010001",
    "1110101011101111",
    "1110100000111001",
    "1110011101001111",
    "1110011111110110",
    "1110100111000011",
    "1110110001001111",
    "1110111101100000",
    "1111001011101000",
    "1111011011101010",
    "1111101101001110",
    "1111111111000101",
    "1111110000101100",
    "1111100100011101",
    "1111011110001001",
    "1111011110100110",
    "1111100101101001",
    "1111110010000011",
    "1111111101111100",
    "1111101100100011",
    "1111011011101101",
    "1111001101000101",
    "1111000010000110",
    "1110111011110111",
    "1110111011000100",
    "1110111111111010",
    "1111001010000100",
    "1111011000110000",
    "1111101010101001",
    "1111111101110001",
    "1111110000000111",
    "1111100001010010",
    "1111010111011101",
    "1111010011011010",
    "1111010100111100",
    "1111011011000110",
    "1111100100011100",
    "1111101111100111",
    "1111111011101101",
    "1111110111100001",
    "1111101001110010",
    "1111011010011101",
    "1111001001010101",
    "1110110111001001",
    "1110100101111100",
    "1110011000011101",
    "1110010001010101",
    "1110010010010100",
    "1110011011100110",
    "1110101011110101",
    "1111000000100110",
    "1111010111010000",
    "1111101101011110",
    "1111111110001100",
    "1111101100111001",
    "1111011111100110",
    "1111010111101101",
    "1111010110110110",
    "1111011110010111",
    "1111101110011011",
    "1111111010100011",
    "1111100000000000",
    "1111000110001110",
    "1110110001010101",
    "1110100100001101",
    "1110011111101001",
    "1110100010101111",
    "1110101011100101",
    "1110111000101101",
    "1111001001100101",
    "1111011110000101",
    "1111110101101010",
    "1111110001001111",
    "1111011001011110",
    "1111000110010110",
    "1110111010101101",
    "1110110111110101",
    "1110111100110011",
    "1111000110111100",
    "1111010010101100",
    "1111011100101101",
    "1111100010101001",
    "1111100011011100",
    "1111011111001010",
    "1111010110101111",
    "1111001011100110",
    "1110111111011010",
    "1110110011110001",
    "1110101010000010",
    "1110100011010000",
    "1110100000001010",
    "1110100001001100",
    "1110100110101010",
    "1110110000100111",
    "1110111110100011",
    "1111001111011001",
    "1111100001100100",
    "1111110011000000",
    "1111111110001100",
    "1111110011100100",
    "1111101101100010",
    "1111101011100101",
    "1111101100011110",
    "1111101110110010",
    "1111110001011000",
    "1111110011101111",
    "1111110101111110",
    "1111111000011100",
    "1111111011010001",
    "1111111101110001",
    "1111111110011111",
    "1111111011100001",
    "1111110011011001",
    "1111100101110110",
    "1111010100001110",
    "1111000001011010",
    "1110110000110000",
    "1110100101010000",
    "1110100000101011",
    "1110100011001000",
    "1110101011100011",
    "1110111000010101",
    "1111001000010011",
    "1111011010110101",
    "1111101111100000",
    "1111111010011001",
    "1111100100010111",
    "1111010000100100",
    "1111000001101001",
    "1110111001100011",
    "1110111001001110",
    "1110111111110110",
    "1111001011010110",
    "1111011001000010",
    "1111100110010010",
    "1111110001000100",
    "1111111000011111",
    "1111111100100100",
    "1111111110001100",
    "1111111110101001",
    "1111111111001011",
    "1111111111010000",
    "1111111100011011",
    "1111111000100010",
    "1111110100001100",
    "1111110000001001",
    "1111101100111101",
    "1111101010110111",
    "1111101001101000",
    "1111101000110000",
    "1111100111110100",
    "1111100110011110",
    "1111100100101001",
    "1111100010010101",
    "1111011111101100",
    "1111011100110011",
    "1111011001110101",
    "1111010111001000",
    "1111010101001101",
    "1111010100110011",
    "1111010110101100",
    "1111011011010100",
    "1111100010101001",
    "1111101100000100",
    "1111110110011111",
    "1111111111010000",
    "1111110110010011",
    "1111101110111110",
    "1111101000111110",
    "1111100011100001",
    "1111011101110101",
    "1111010111100111",
    "1111010001001100",
    "1111001011100001",
    "1111000111110111",
    "1111000111010011",
    "1111001010010001",
    "1111010000011111",
    "1111011000111100",
    "1111100010001000",
    "1111101010010001",
    "1111101111101000",
    "1111110000110011",
    "1111101101000010",
    "1111100100010000",
    "1111010111001000",
    "1111000110110111",
    "1110110101010111",
    "1110100100101001",
    "1110010110110001",
    "1110001101000111",
    "1110001000010011",
    "1110000111110101",
    "1110001010011110",
    "1110001110100110",
    "1110010010111001",
    "1110010111101101",
    "1110011110101011",
    "1110101001100000",
    "1110111000101000",
    "1111001010011000",
    "1111011011011000",
    "1111100111100010",
    "1111101011101000",
    "1111100110101001",
    "1111011010011110",
    "1111001010111101",
    "1110111100011110",
    "1110110010010010",
    "1110101101101110",
    "1110101110010110",
    "1110110010010010",
    "1110110111001000",
    "1110111010110101",
    "1110111100001010",
    "1110111010110111",
    "1110110111011111",
    "1110110011010111",
    "1110110000010100",
    "1110110000011001",
    "1110110101111110",
    "1111000011010000",
    "1111011001001100",
    "1111110110011110",
    "1111101000100111",
    "1111001001011011",
    "1110110001001111",
    "1110100011111011",
    "1110100010101001",
    "1110101011101010",
    "1110111010111101",
    "1111001011111100",
    "1111011010101111",
    "1111100101010011",
    "1111101011010100",
    "1111101111010101",
    "1111110110011011",
    "1111111010111111",
    "1111100011111011",
    "1111000111010101",
    "1110101011011001",
    "1110010110101010",
    "1110001101110101",
    "1110010010100010",
    "1110100001110000",
    "1110110101101111",
    "1111001000110000",
    "1111010110100111",
    "1111011101111111",
    "1111011111111010",
    "1111011110011111",
    "1111011101001111",
    "1111011111101000",
    "1111100111010111",
    "1111110100000011",
    "1111111100111011",
    "1111101111101011",
    "1111100111011100",
    "1111100101101110",
    "1111101001101001",
    "1111110000000110",
    "1111110100100010",
    "1111110010011011",
    "1111100110111111",
    "1111010010110110",
    "1110111001110000",
    "1110100001000000",
    "1110001101100100",
    "1110000010100100",
    "1110000000011100",
    "1110000101101111",
    "1110001111111111",
    "1110011101001001",
    "1110101100100000",
    "1110111110011111",
    "1111010011100111",
    "1111101011011011",
    "1111111011110000",
    "1111100100100000",
    "1111010001011010",
    "1111000100011101",
    "1110111110000111",
    "1110111101001010",
    "1110111111011110",
    "1111000010111001",
    "1111000110010101",
    "1111001010000110",
    "1111001111001100",
    "1111010110011011",
    "1111011111110110",
    "1111101010010101",
    "1111110100010000",
    "1111111100000000",
    "1111111111101000",
    "1111111111000101",
    "1111111110010001",
    "1111111001110011",
    "1111110100110010",
    "1111110000001100",
    "1111101100100100",
    "1111101010000100",
    "1111101000100111",
    "1111101000000010",
    "1111101000010001",
    "1111101001100000",
    "1111101100001010",
    "1111110000010010",
    "1111110101111101",
    "1111111101101111",
    "1111110110111011",
    "1111100110111001",
    "1111010010001010",
    "1110111010110100",
    "1110100100011101",
    "1110010011000000",
    "1110001001100000",
    "1110001001000111",
    "1110010001000000",
    "1110011111000111",
    "1110110001011110",
    "1111000110100010",
    "1111011101000100",
    "1111110011010000",
    "1111111001011000",
    "1111101011101111",
    "1111100110010011",
    "1111101010100100",
    "1111111000100111",
    "1111110000010000",
    "1111010001111000",
    "1110101110111010",
    "1110001010110111",
    "1101101001101111",
    "1101001111010100",
    "1100111110011100",
    "1100111000101100",
    "1100111101100000",
    "1101001010001110",
    "1101011011000100",
    "1101101100000111",
    "1101111010100011",
    "1110000101010011",
    "1110001100111111",
    "1110010100101010",
    "1110100001001101",
    "1110110110010011",
    "1111010100110100",
    "1111111001110010",
    "1111100000101100",
    "1111000001010101",
    "1110101101010111",
    "1110100111001000",
    "1110101100110010",
    "1110111001101010",
    "1111001000001011",
    "1111010011110110",
    "1111011010100110",
    "1111011100101010",
    "1111011011100110",
    "1111011011000100",
    "1111011111101100",
    "1111101100101110",
    "1111111101000011",
    "1111100000010111",
    "1111000010010111",
    "1110101000101101",
    "1110010111110101",
    "1110010001110100",
    "1110010101001101",
    "1110011110010100",
    "1110101000100111",
    "1110110000011100",
    "1110110100011111",
    "1110110101011101",
    "1110110100111110",
    "1110110100110110",
    "1110110101111001",
    "1110110111101101",
    "1110111001010001",
    "1110111001010110",
    "1110110111011000",
    "1110110100001011",
    "1110110001011110",
    "1110110001001111",
    "1110110101010111",
    "1110111111010010",
    "1111010000000010",
    "1111100111101101",
    "1111111011010001",
    "1111011100001110",
    "1110111111010001",
    "1110101000010011",
    "1110011001110101",
    "1110010100100010",
    "1110010111001011",
    "1110011111100001",
    "1110101011100101",
    "1110111010100110",
    "1111001100110111",
    "1111100010100110",
    "1111111011000010",
    "1111101011111110",
    "1111010101011111",
    "1111000100001110",
    "1110111001110111",
    "1110110110010110",
    "1110111000010110",
    "1110111110001100",
    "1111000110100101",
    "1111010001011110",
    "1111011111010100",
    "1111110000010110",
    "1111111100010101",
    "1111101001001100",
    "1111011001011000",
    "1111001111110110",
    "1111001110010001",
    "1111010100100000",
    "1111100000101001",
    "1111101111100011",
    "1111111101111111",
    "1111110110010100",
    "1111101110011000",
    "1111101010001111",
    "1111101001010111",
    "1111101011010110",
    "1111101111110101",
    "1111110110101101",
    "1111111111111110",
    "1111110100011010",
    "1111100110111100",
    "1111011000001011",
    "1111001000110111",
    "1110111001111010",
    "1110101100011100",
    "1110100001101110",
    "1110011010111100",
    "1110011000111001",
    "1110011011110101",
    "1110100011011010",
    "1110101110011110",
    "1110111011110111",
    "1111001011110011",
    "1111011111101000",
    "1111111000010011",
    "1111101011000000",
    "1111001101111000",
    "1110110101100000",
    "1110100111000100",
    "1110100101110110",
    "1110110001101110",
    "1111000111010011",
    "1111100010000011",
    "1111111110101001",
    "1111100100000000",
    "1111000101100010",
    "1110100101101111",
    "1110000110000011",
    "1101101001100101",
    "1101010100100111",
    "1101001011000001",
    "1101001110100100",
    "1101011110111101",
    "1101111001111111",
    "1110011100010011",
    "1111000001111101",
    "1111100111000101",
    "1111110111111010",
    "1111011110000010",
    "1111001101010111",
    "1111000110100000",
    "1111001000001001",
    "1111001111011100",
    "1111011000111010",
    "1111100001101011",
    "1111101000001100",
    "1111101100011000",
    "1111101111000010",
    "1111110001010011",
    "1111110011110011",
    "1111110110011110",
    "1111111000111100",
    "1111111011000110",
    "1111111101011010",
    "1111111111001110",
    "1111111010010011",
    "1111110011111100",
    "1111101101001110",
    "1111100111110100",
    "1111100101010011",
    "1111100110100010",
    "1111101011000011",
    "1111110001000101",
    "1111110110001011",
    "1111111000000010",
    "1111110101010000",
    "1111101101101110",
    "1111100010100111",
    "1111010101101100",
    "1111001000110010",
    "1110111101001110",
    "1110110011101100",
    "1110101100011100",
    "1110100111100011",
    "1110100101011000",
    "1110100110100100",
    "1110101011101000",
    "1110110100101001",
    "1111000001010000",
    "1111010000110101",
    "1111100010100001",
    "1111110101011010",
    "1111110111011100",
    "1111100101010010",
    "1111010101001101",
    "1111001000011010",
    "1110111111100110",
    "1110111011000111",
    "1110111010101111",
    "1110111101110111",
    "1111000011110110",
    "1111001100010100",
    "1111010111000001",
    "1111100011111011",
    "1111110010101000",
    "1111111101100111",
    "1111101110010101",
    "1111100001100010",
    "1111011001010110",
    "1111010111011011",
    "1111011100010110",
    "1111100111001101",
    "1111110101101001",
    "1111111011011101",
    "1111101111011101",
    "1111101000110101",
    "1111101000110111",
    "1111101111101010",
    "1111111100011110",
    "1111110010000100",
    "1111011101110101",
    "1111001000111111",
    "1110110101110100",
    "1110100110010110",
    "1110011100000001",
    "1110010111010011",
    "1110010111101010",
    "1110011011110010",
    "1110100001111000",
    "1110101000110000",
    "1110110000100100",
    "1110111010111100",
    "1111001001111111",
    "1111011110110110",
    "1111111000110011",
    "1111101011000011",
    "1111010001010010",
    "1110111110011001",
    "1110110101010011",
    "1110110110011011",
    "1110111111110110",
    "1111001110011100",
    "1111011111000101",
    "1111101111110000",
    "1111111111110000",
    "1111110000100010",
    "1111100000010111",
    "1111001111010110",
    "1110111110000010",
    "1110101110000100",
    "1110100001011100",
    "1110011010000001",
    "1110011000101010",
    "1110011101000111",
    "1110100110000011",
    "1110110001100100",
    "1110111101101101",
    "1111001000111111",
    "1111010011101110",
    "1111011111110110",
    "1111101111110100",
    "1111111011010011",
    "1111100011000000",
    "1111001011001001",
    "1110111000101101",
    "1110110000010100",
    "1110110100011000",
    "1111000011111011",
    "1111011010111101",
    "1111110100001001",
    "1111110101111011",
    "1111100111100001",
    "1111100011001000",
    "1111101001101010",
    "1111111001111110",
    "1111101110100100",
    "1111010011100111",
    "1110111001010001",
    "1110100011010111",
    "1110010100100010",
    "1110001101111111",
    "1110001111001000",
    "1110010101111100",
    "1110011111011010",
    "1110101000110100",
    "1110110000100110",
    "1110110111100111",
    "1111000000011001",
    "1111001101101000",
    "1111100000001000",
    "1111110110010110",
    "1111110011010110",
    "1111100001011110",
    "1111010111100000",
    "1111010110110010",
    "1111011101101000",
    "1111101000011010",
    "1111110011001110",
    "1111111011010010",
    "1111111111110101",
    "1111111110001001",
    "1111111100111100",
    "1111111010101110",
    "1111110110100110",
    "1111110000011111",
    "1111101001000000",
    "1111100000111101",
    "1111011001010110",
    "1111010011000101",
    "1111001110111000",
    "1111001101010100",
    "1111001110101001",
    "1111010010100111",
    "1111011000011101",
    "1111011111011110",
    "1111100111011000",
    "1111110000011111",
    "1111111011011111",
    "1111110111000101",
    "1111100111100111",
    "1111010111010001",
    "1111001000000011",
    "1110111011111111",
    "1110110100100100",
    "1110110010001011",
    "1110110100001011",
    "1110111001000010",
    "1110111111011100",
    "1111000111000001",
    "1111010000110000",
    "1111011110001001",
    "1111110000000100",
    "1111111010001001",
    "1111100011001011",
    "1111001110110000",
    "1111000000101110",
    "1110111011011000",
    "1110111110111011",
    "1111001001100010",
    "1111011000001011",
    "1111100111101000",
    "1111110101010100",
    "1111111111100001",
    "1111111010101011",
    "1111111001100111",
    "1111111101001110",
    "1111111010100110",
    "1111101110100110",
    "1111100000000011",
    "1111010000110011",
    "1111000010110011",
    "1110110111110010",
    "1110110000101100",
    "1110101101110011",
    "1110101110100100",
    "1110110010000110",
    "1110110111011011",
    "1110111101110000",
    "1111000100101001",
    "1111001100100001",
    "1111010110101101",
    "1111100100111001",
    "1111111000010001",
    "1111101111011010",
    "1111010100010111",
    "1110111010001111",
    "1110100101010000",
    "1110011000101101",
    "1110010101111011",
    "1110011011111101",
    "1110101000001011",
    "1110110111001110",
    "1111000101111110",
    "1111010010001101",
    "1111011010110000",
    "1111011111011001",
    "1111100000011111",
    "1111011110011001",
    "1111011001100101",
    "1111010010100001",
    "1111001010000001",
    "1111000001001101",
    "1110111001100011",
    "1110110100010101",
    "1110110010010000",
    "1110110011010010",
    "1110110110101000",
    "1110111011001110",
    "1110111111110110",
    "1111000011110110",
    "1111000111110111",
    "1111001110100011",
    "1111011011100011",
    "1111110001010000",
    "1111110000111000",
    "1111001111000000",
    "1110101111001010",
    "1110010111100111",
    "1110001100101101",
    "1110001111011001",
    "1110011101010110",
    "1110110010110100",
    "1111001100000010",
    "1111100110000100",
    "1111111110101111",
    "1111101100000110",
    "1111011100110111",
    "1111010101110100",
    "1111011001001001",
    "1111101000000001",
    "1111111110010110",
    "1111011101000010",
    "1110111000110100",
    "1110010111001101",
    "1101111101000100",
    "1101101101011001",
    "1101101000111010",
    "1101101110011100",
    "1101111100001001",
    "1110010000000111",
    "1110101000111001",
    "1111000101000001",
    "1111100010101100",
    "1111111111101011",
    "1111100110100000",
    "1111010010000010",
    "1111000011111001",
    "1110111011101000",
    "1110110111101100",
    "1110110110011000",
    "1110110110011101",
    "1110110111101010",
    "1110111010011011",
    "1110111111011110",
    "1111000110111110",
    "1111010000001010",
    "1111011001010001",
    "1111100000100100",
    "1111100100101111",
    "1111100101110110",
    "1111100110101010",
    "1111101011110110",
    "1111111000110101",
    "1111110001111100",
    "1111010111110001",
    "1110111101111111",
    "1110101001111010",
    "1110011111001101",
    "1110011110001100",
    "1110100011011100",
    "1110101010000110",
    "1110101110001001",
    "1110101110010100",
    "1110101100111000",
    "1110101101101011",
    "1110110100000001",
    "1111000001010000",
    "1111010011100010",
    "1111100110011100",
    "1111110100110111",
    "1111111010011100",
    "1111110101001101",
    "1111100110011010",
    "1111010001100100",
    "1110111010111100",
    "1110100110001110",
    "1110010110010010",
    "1110001101000000",
    "1110001011010011",
    "1110010000100110",
    "1110011100010011",
    "1110101101111111",
    "1111000101001101",
    "1111100000110110",
    "1111111110100011",
    "1111100101001001",
    "1111001101110011",
    "1110111101110111",
    "1110110110010110",
    "1110110110100101",
    "1110111101001010",
    "1111001000110100",
    "1111011001000110",
    "1111101101110111",
    "1111111001100100",
    "1111011111010111",
    "1111000110101101",
    "1110110011001011",
    "1110100111011011",
    "1110100100010010",
    "1110101000101101",
    "1110110010011101",
    "1110111111000111",
    "1111001100111010",
    "1111011011011011",
    "1111101010111100",
    "1111111011110000",
    "1111110010110101",
    "1111100011000000",
    "1111010111100000",
    "1111010010011101",
    "1111010100110100",
    "1111011110000111",
    "1111101100110110",
    "1111111110111000",
    "1111101110000111",
    "1111011100010001",
    "1111001101001001",
    "1111000010000011",
    "1110111100001001",
    "1110111100010001",
    "1111000010100110",
    "1111001110101101",
    "1111011111011110",
    "1111110011100000",
    "1111110110100101",
    "1111100000001100",
    "1111001010100101",
    "1110110110111110",
    "1110100110100000",
    "1110011010011101",
    "1110010011111000",
    "1110010011011111",
    "1110011001010001",
    "1110100101001110",
    "1110110111110101",
    "1111010001000000",
    "1111101111001000",
    "1111110001011001",
    "1111010101110010",
    "1111000010110100",
    "1110111011110101",
    "1111000001101100",
    "1111010010101100",
    "1111101011101100",
    "1111110110011011",
    "1111010110100000",
    "1110110110111111",
    "1110011010011001",
    "1110000011101001",
    "1101110101100111",
    "1101110010100001",
    "1101111011100101",
    "1110010000101100",
    "1110110000011111",
    "1111010111111100",
    "1111111101101101",
    "1111010110010010",
    "1110110110111011",
    "1110100011000000",
    "1110011011100101",
    "1110011111001111",
    "1110101010110101",
    "1110111010011011",
    "1111001010001100",
    "1111010111101101",
    "1111100001111000",
    "1111101001000100",
    "1111101110101101",
    "1111110100111110",
    "1111111110001011",
    "1111110011111010",
    "1111100000111000",
    "1111001001110111",
    "1110110001100110",
    "1110011011101111",
    "1110001011101111",
    "1110000011110100",
    "1110000100001101",
    "1110001010110111",
    "1110010100010010",
    "1110011101000100",
    "1110100100001000",
    "1110101100001010",
    "1110111001001011",
    "1111001101100011",
    "1111101000000110",
    "1111111011110111",
    "1111100100100100",
    "1111010111001011",
    "1111010110001011",
    "1111011111100001",
    "1111101101100111",
    "1111111010010100",
    "1111111110101101",
    "1111111110100110",
    "1111111100100111",
    "1111110110011001",
    "1111110010110001",
    "1111110100110111",
    "1111111101001010",
    "1111110110100100",
    "1111101010100100",
    "1111100011100010",
    "1111100100110011",
    "1111101111010011",
    "1111111110011001",
    "1111100111110111",
    "1111010001011100",
    "1110111111100001",
    "1110110101010101",
    "1110110100000000",
    "1110111010110010",
    "1111001000001001",
    "1111011010110000",
    "1111110001101010",
    "1111110100001010",
    "1111011000101000",
    "1110111110100001",
    "1110101000111110",
    "1110011011000111",
    "1110010110111100",
    "1110011100100110",
    "1110101010100011",
    "1110111110011110",
    "1111010101111100",
    "1111101110110001",
    "1111111001001101",
    "1111100100010111",
    "1111010100101001",
    "1111001011101101",
    "1111001010100011",
    "1111010001101001",
    "1111100000101110",
    "1111110110100111",
    "1111101110110111",
    "1111010010100001",
    "1110110111001101",
    "1110011111001010",
    "1110001011110101",
    "1101111101110000",
    "1101110100110011",
    "1101110000010100",
    "1101101111111011",
    "1101110100000110",
    "1101111110010110",
    "1110010000000010",
    "1110101001000100",
    "1111000111001000",
    "1111100101111001",
    "1111111111111001",
    "1111101111010100",
    "1111101011011011",
    "1111110100010110",
    "1111111000100110",
    "1111011111110101",
    "1111000101111100",
    "1110101111000000",
    "1110011101110011",
    "1110010011110001",
    "1110010000110101",
    "1110010011111100",
    "1110011011101010",
    "1110100110110010",
    "1110110100101100",
    "1111000101100101",
    "1111011010010110",
    "1111110100000001",
    "1111101101010011",
    "1111001011100000",
    "1110101010011001",
    "1110001110111000",
    "1101111101010110",
    "1101111000001011",
    "1101111110110011",
    "1110001110000100",
    "1110100001110100",
    "1110110111101101",
    "1111010000001100",
    "1111101100111010",
    "1111110001011101",
    "1111001100111100",
    "1110101010001110",
    "1110001111011001",
    "1110000001101100",
    "1110000011011010",
    "1110010010011101",
    "1110101001100101",
    "1111000011010011",
    "1111011100101010",
    "1111110101100110",
    "1111110000011100",
    "1111010101000000",
    "1110111001100111",
    "1110100010001010",
    "1110010011010101",
    "1110010000011111",
    "1110011001011110",
    "1110101010100010",
    "1110111101101101",
    "1111001101001001",
    "1111010101001101",
    "1111010101010101",
    "1111001111011001",
    "1111000110101010",
    "1110111110101011",
    "1110111010011000",
    "1110111011110101",
    "1111000011101111",
    "1111010001100010",
    "1111100011011000",
    "1111110110101000",
    "1111110111100100",
    "1111101001110110",
    "1111100001110000",
    "1111011111010001",
    "1111100001000111",
    "1111100101010111",
    "1111101010011001",
    "1111101111011100",
    "1111110100011001",
    "1111111001011001",
    "1111111110010111",
    "1111111101010000",
    "1111111010101101",
    "1111111011011101",
    "1111111111011010",
    "1111110110000011",
    "1111101001111110",
    "1111011101101000",
    "1111010011011111",
    "1111001101010010",
    "1111001011100110",
    "1111001101110101",
    "1111010010110110",
    "1111011001100011",
    "1111100001011100",
    "1111101010110101",
    "1111110110011101",
    "1111111011001100",
    "1111101010010011",
    "1111010111100111",
    "1111000100011100",
    "1110110010011101",
    "1110100011101110",
    "1110011010000111",
    "1110010110111100",
    "1110011010101011",
    "1110100101000110",
    "1110110101001011",
    "1111001001001001",
    "1111011110011110",
    "1111110010010001",
    "1111111110010010",
    "1111110101110001",
    "1111110101101101",
    "1111111110010110",
    "1111110001101100",
    "1111011101010111",
    "1111001000010101",
    "1110110110001110",
    "1110101001110010",
    "1110100100011101",
    "1110100110010000",
    "1110101110010110",
    "1110111011001111",
    "1111001011010100",
    "1111011100111101",
    "1111101110011011",
    "1111111101111111",
    "1111110101110000",
    "1111101101110110",
    "1111101010011001",
    "1111101010111101",
    "1111101110111101",
    "1111110110000111",
    "1111111111011000",
    "1111110001001110",
    "1111011111100011",
    "1111001011011011",
    "1110110111000100",
    "1110100101010011",
    "1110011000111001",
    "1110010011110001",
    "1110010110101111",
    "1110100001010100",
    "1110110010001000",
    "1111000111011011",
    "1111011111011100",
    "1111111000011001",
    "1111101111010110",
    "1111011001100010",
    "1111000111101010",
    "1110111010111100",
    "1110110011111110",
    "1110110010011101",
    "1110110101100100",
    "1110111100000100",
    "1111000100101100",
    "1111001110011100",
    "1111011000101000",
    "1111100010101100",
    "1111101100011111",
    "1111110110101101",
    "1111111101000010",
    "1111101101001001",
    "1111011001000110",
    "1111000010010111",
    "1110101100001010",
    "1110011010011000",
    "1110010000001111",
    "1110001110111111",
    "1110010101001110",
    "1110011111101110",
    "1110101010101000",
    "1110110010111001",
    "1110110111001001",
    "1110110111100111",
    "1110110101011101",
    "1110110010001010",
    "1110101110110011",
    "1110101011111101",
    "1110101001101111",
    "1110101000010000",
    "1110100111111111",
    "1110101010011110",
    "1110110001111101",
    "1111000000100110",
    "1111010111001101",
    "1111110100100001",
    "1111101010110010",
    "1111001011011000",
    "1110110001101100",
    "1110100000111011",
    "1110011001111001",
    "1110011011000001",
    "1110100001001111",
    "1110101001010000",
    "1110110000011100",
    "1110110101011011",
    "1110110111110010",
    "1110110111101000",
    "1110110101100100",
    "1110110010010010",
    "1110101110110110",
    "1110101100010111",
    "1110101011111101",
    "1110101110010111",
    "1110110100000110",
    "1110111110001101",
    "1111001110011011",
    "1111100101101110",
    "1111111100101100",
    "1111011100001010",
    "1110111101101110",
    "1110100110100111",
    "1110011010110101",
    "1110011011100011",
    "1110100110011111",
    "1110110110111001",
    "1111000111101101",
    "1111010101000101",
    "1111011101011100",
    "1111100001011001",
    "1111100010111011",
    "1111100101000110",
    "1111101010110000",
    "1111110101011010",
    "1111111011011011",
    "1111101010011011",
    "1111011011011011",
    "1111010010001111",
    "1111010001100010",
    "1111011010001111",
    "1111101011000011",
    "1111111111001000",
    "1111101000100101",
    "1111010101010011",
    "1111001000010000",
    "1111000010111101",
    "1111000101110001",
    "1111010000010001",
    "1111100001001010",
    "1111110110011100",
    "1111110010101111",
    "1111011101100001",
    "1111001100101000",
    "1111000001111011",
    "1110111101111111",
    "1110111111110001",
    "1111000101001000",
    "1111001011101010",
    "1111010001101110",
    "1111010110101010",
    "1111011010110010",
    "1111011110101001",
    "1111100010101100",
    "1111100110110000",
    "1111101001110101",
    "1111101010011101",
    "1111100111001110",
    "1111011111100011",
    "1111010100000000",
    "1111000110001011",
    "1110111000001011",
    "1110101011101011",
    "1110100001111001",
    "1110011011011101",
    "1110011000100111",
    "1110011001101000",
    "1110011110111010",
    "1110101001000111",
    "1110111000110111",
    "1111001110001010",
    "1111100111111000",
    "1111111100000011",
    "1111100000100001",
    "1111001000001011",
    "1110110101001000",
    "1110101000011011",
    "1110100010000010",
    "1110100000111110",
    "1110100011111000",
    "1110101001010001",
    "1110101111101100",
    "1110110101111100",
    "1110111010111010",
    "1110111110000010",
    "1110111111010010",
    "1110111111101100",
    "1111000001100111",
    "1111001000000110",
    "1111010101100000",
    "1111101010010001",
    "1111111011110011",
    "1111100001000101",
    "1111001010011001",
    "1110111011101111",
    "1110110110101111",
    "1110111010001001",
    "1111000010111001",
    "1111001101001111",
    "1111010110010010",
    "1111011100001010",
    "1111011110000101",
    "1111011011110111",
    "1111010101101001",
    "1111001011111111",
    "1110111111111011",
    "1110110011010101",
    "1110101000110111",
    "1110100011100001",
    "1110100110010000",
    "1110110011001101",
    "1111001010100110",
    "1111101010001110",
    "1111110010010001",
    "1111010000001101",
    "1110110100010011",
    "1110100001110001",
    "1110011001010110",
    "1110011001100011",
    "1110011111001111",
    "1110100110101111",
    "1110101101010010",
    "1110110001100010",
    "1110110011011111",
    "1110110100001000",
    "1110110100111011",
    "1110110111000110",
    "1110111011011011",
    "1111000001111110",
    "1111001010110101",
    "1111010111000110",
    "1111101000100101",
    "1111111111011111",
    "1111100001111000",
    "1111000001100111",
    "1110100011011000",
    "1110001011110111",
    "1101111110011100",
    "1101111100000010",
    "1110000010011100",
    "1110001101101101",
    "1110011001100010",
    "1110100011010000",
    "1110101011010011",
    "1110110100100010",
    "1111000010010000",
    "1111010110001110",
    "1111101111010000",
    "1111110110100001",
    "1111100000011010",
    "1111010011001011",
    "1111010001010101",
    "1111011010010001",
    "1111101011001000",
    "1111111111100110",
    "1111101001001011",
    "1111010011110100",
    "1111000001010100",
    "1110110011000000",
    "1110101001101101",
    "1110100101110100",
    "1110100111011010",
    "1110101110001111",
    "1110111010000010",
    "1111001010010110",
    "1111011110000010",
    "1111110011010010",
    "1111111000010001",
    "1111100111100010",
    "1111011101001111",
    "1111011011101000",
    "1111100011100110",
    "1111110100011100",
    "1111110100001100",
    "1111011001111111",
    "1111000001000011",
    "1110101100110010",
    "1110011111010110",
    "1110011001011011",
    "1110011010011110",
    "1110100000111011",
    "1110101010110111",
    "1110110110100100",
    "1111000011001111",
    "1111010001101100",
    "1111100011110001",
    "1111111011000110",
    "1111101000010011",
    "1111001000110101",
    "1110101010101111",
    "1110010010100100",
    "1110000011111001",
    "1101111111111000",
    "1110000101001110",
    "1110010001001000",
    "1110100000011111",
    "1110110001000011",
    "1111000001110001",
    "1111010010010101",
    "1111100010100111",
    "1111110010001010",
    "1111111111111100",
    "1111110101000001",
    "1111101110000001",
    "1111101011001001",
    "1111101011110011",
    "1111101110101011",
    "1111110010010101",
    "1111110101101011",
    "1111111000010010",
    "1111111010001000",
    "1111111011010110",
    "1111111100000001",
    "1111111100001110",
    "1111111100000100",
    "1111111011101110",
    "1111111011010001",
    "1111111010100100",
    "1111111001010010",
    "1111110110111010",
    "1111110011000111",
    "1111101110000011",
    "1111101000011110",
    "1111100011101001",
    "1111100001000101",
    "1111100010011100",
    "1111101001010011",
    "1111110110111000",
    "1111110100100101",
    "1111011010110000",
    "1110111110111111",
    "1110100101100100",
    "1110010010100001",
    "1110001000101000",
    "1110001000101010",
    "1110010001011111",
    "1110100001001000",
    "1110110110001110",
    "1111010000010001",
    "1111101110110111",
    "1111101111011100",
    "1111001101110011",
    "1110110000011100",
    "1110011011011110",
    "1110010001110000",
    "1110010011111011",
    "1110100000111110",
    "1110110110111011",
    "1111010011010111",
    "1111110011100101",
    "1111101011100010",
    "1111001101010100",
    "1110110100101111",
    "1110100100001011",
    "1110011100100110",
    "1110011101000111",
    "1110100011001011",
    "1110101011101000",
    "1110110100001000",
    "1110111011101111",
    "1111000011001101",
    "1111001100101000",
    "1111011010001111",
    "1111101101010000",
    "1111111011001001",
    "1111100001110100",
    "1111001010100101",
    "1110111000110010",
    "1110101110010111",
    "1110101011010100",
    "1110101110001111",
    "1110110100110100",
    "1110111100111000",
    "1111000101010101",
    "1111001110110011",
    "1111011011000001",
    "1111101011001000",
    "1111111110110000",
    "1111101100101101",
    "1111011011100000",
    "1111010001110000",
    "1111010010001101",
    "1111011101010100",
    "1111110001010110",
    "1111110100101000",
    "1111011000011000",
    "1110111101011100",
    "1110100110111110",
    "1110010111011111",
    "1110010000100100",
    "1110010010100100",
    "1110011100011011",
    "1110101011101111",
    "1110111101100100",
    "1111001111001010",
    "1111011110010111",
    "1111101001111001",
    "1111110001100001",
    "1111110110001011",
    "1111111010011111",
    "1111111110001100",
    "1111110001110010",
    "1111100000011111",
    "1111001101001010",
    "1110111100011100",
    "1110110011000011",
    "1110110100010101",
    "1111000000111011",
    "1111010110001000",
    "1111101111001110",
    "1111111000110001",
    "1111100101111100",
    "1111011010001110",
    "1111010101110010",
    "1111010111110001",
    "1111011110011011",
    "1111101000010011",
    "1111110100001100",
    "1111111110111010",
    "1111110010000010",
    "1111100110000011",
    "1111011011111101",
    "1111010100100101",
    "1111010000010101",
    "1111001111010110",
    "1111010001011110",
    "1111010110101100",
    "1111011110101001",
    "1111101000011111",
    "1111110011001000",
    "1111111101011011",
    "1111111001100001",
    "1111110010010101",
    "1111101101010000",
    "1111101010100110",
    "1111101010111100",
    "1111101111000111",
    "1111110111110110",
    "1111111010110110",
    "1111101010000110",
    "1111010111110100",
    "1111000110100010",
    "1110111000101000",
    "1110110000000011",
    "1110101110000000",
    "1110110010111101",
    "1110111110100011",
    "1111001111110110",
    "1111100101010101",
    "1111111101000001",
    "1111101011011101",
    "1111010110100101",
    "1111000110011011",
    "1110111100011011",
    "1110111001000010",
    "1110111011110010",
    "1111000011001111",
    "1111001101100110",
    "1111011001001110",
    "1111100110001000",
    "1111110110001100",
    "1111110100010111",
    "1111011001000010",
    "1110111010000001",
    "1110011011110011",
    "1110000011100111",
    "1101110101101001",
    "1101110011010111",
    "1101111010110101",
    "1110000111110001",
    "1110010101100100",
    "1110100001100010",
    "1110101100110011",
    "1110111011000100",
    "1111001111100100",
    "1111101010111100",
    "1111110110001110",
    "1111011010100101",
    "1111001001011000",
    "1111001000100010",
    "1111011001111111",
    "1111111010011010",
    "1111011101010111",
    "1110110101110111",
    "1110010110001110",
    "1110000010011101",
    "1101111100000010",
    "1110000010000011",
    "1110010001101110",
    "1110101000000110",
    "1111000010011101",
    "1111011110101000",
    "1111111010101000",
    "1111101011011111",
    "1111010110000000",
    "1111000110011111",
    "1110111101010110",
    "1110111001110100",
    "1110111010001110",
    "1110111100111101",
    "1111000000101011",
    "1111000100011111",
    "1111001000000110",
    "1111001011100101",
    "1111001111001100",
    "1111010011001111",
    "1111010111111001",
    "1111011101110010",
    "1111100110001001",
    "1111110010100000",
    "1111111100100000",
    "1111100111111001",
    "1111010010100001",
    "1111000000010100",
    "1110110100111011",
    "1110110010011100",
    "1110111000011101",
    "1111000100000101",
    "1111010001010101",
    "1111011100101011",
    "1111100100000001",
    "1111100110111111",
    "1111100110010011",
    "1111100011001010",
    "1111011111001101",
    "1111011100100110",
    "1111011101101011",
    "1111100100001000",
    "1111110000011000",
    "1111111110110100",
    "1111101100010001",
    "1111011011101101",
    "1111010000110110",
    "1111001110001010",
    "1111010011100100",
    "1111011110011111",
    "1111101010111011",
    "1111110100110010",
    "1111111001001000",
    "1111110110110000",
    "1111101110010011",
    "1111100001111000",
    "1111010100000001",
    "1111000110111110",
    "1110111100001110",
    "1110110100100101",
    "1110110000011001",
    "1110101111110101",
    "1110110011000001",
    "1110111010001100",
    "1111000101011010",
    "1111010100011010",
    "1111100110010101",
    "1111111001011111",
    "1111110100001101",
    "1111100101000000",
    "1111011010010100",
    "1111010100101110",
    "1111010011100100",
    "1111010101100100",
    "1111011001000100",
    "1111011100111111",
    "1111100000111001",
    "1111100101001110",
    "1111101010110011",
    "1111110010001000",
    "1111111010110111",
    "1111111100011011",
    "1111110110000001",
    "1111110011111100",
    "1111110111011110",
    "1111111111010110",
    "1111110001110111",
    "1111100010001101",
    "1111010010101110",
    "1111000101010011",
    "1110111011001111",
    "1110110101001101",
    "1110110011010111",
    "1110110101101111",
    "1110111100010001",
    "1111000111000001",
    "1111010101111100",
    "1111101000110000",
    "1111111110101101",
    "1111101001011111",
    "1111010001110100",
    "1110111100011011",
    "1110101011011001",
    "1110100000000111",
    "1110011011000111",
    "1110011011111010",
    "1110100001010000",
    "1110101001100000",
    "1110110011010000",
    "1110111110010110",
    "1111001011111100",
    "1111011101011110",
    "1111110011010010",
    "1111110100001100",
    "1111011100100110",
    "1111001010010001",
    "1111000001000000",
    "1111000010100111",
    "1111001110001001",
    "1111100000010100",
    "1111110101000000",
    "1111110111101100",
    "1111101000101110",
    "1111011111101000",
    "1111011101001010",
    "1111100001011111",
    "1111101100001111",
    "1111111100100100",
    "1111101111011100",
    "1111011010100110",
    "1111000111111010",
    "1110111001110111",
    "1110110001110011",
    "1110101111100001",
    "1110110001100001",
    "1110110101110001",
    "1110111010101000",
    "1110111111100011",
    "1111000100101001",
    "1111001010011001",
    "1111010001001010",
    "1111011000110100",
    "1111100000110000",
    "1111101000001100",
    "1111101110100000",
    "1111110011101011",
    "1111111000100011",
    "1111111110101100",
    "1111111000000101",
    "1111101010101011",
    "1111011001010001",
    "1111000101100101",
    "1110110010011001",
    "1110100010011100",
    "1110010111110100",
    "1110010011001000",
    "1110010011100001",
    "1110010111000001",
    "1110011011010001",
    "1110011110010001",
    "1110011110110011",
    "1110011100110010",
    "1110011001011101",
    "1110010111001110",
    "1110011000100000",
    "1110011110100100",
    "1110101000101111",
    "1110110100010101",
    "1110111101100110",
    "1111000000110110",
    "1110111011110101",
    "1110101110101101",
    "1110011100000101",
    "1110001000010000",
    "1101110111101100",
    "1101101101101110",
    "1101101011110011",
    "1101110001100100",
    "1101111101100001",
    "1110001110011011",
    "1110100100000001",
    "1110111110011001",
    "1111011100111111",
    "1111111101101001",
    "1111100011001010",
    "1111001001100111",
    "1110111000111010",
    "1110110010000011",
    "1110110011100010",
    "1110111010001001",
    "1111000010011001",
    "1111001001111100",
    "1111010000001000",
    "1111010101110001",
    "1111011100000111",
    "1111100100000011",
    "1111101101010001",
    "1111110110010100",
    "1111111101001111",
    "1111111111101011",
    "1111111110101001",
    "1111111000110011",
    "1111110000001000",
    "1111100110011110",
    "1111011101101101",
    "1111010111011000",
    "1111010100110110",
    "1111010111010110",
    "1111011111111000",
    "1111101110110001",
    "1111111100100011",
    "1111100100000000",
    "1111001010000100",
    "1110110001100001",
    "1110011100101110",
    "1110001101100000",
    "1110000100101110",
    "1110000010011101",
    "1110000110001101",
    "1110001110111010",
    "1110011011100001",
    "1110101011000001",
    "1110111100101101",
    "1111010000000111",
    "1111100100110011",
    "1111111001111001",
    "1111110001110111",
    "1111100000001100",
    "1111010010101011",
    "1111001010100000",
    "1111001000000001",
    "1111001010100010",
    "1111010000100111",
    "1111011000101101",
    "1111100001100111",
    "1111101010111101",
    "1111110100111010",
    "1111111111110011",
    "1111110100101100",
    "1111101001110010",
    "1111100001010100",
    "1111011101000101",
    "1111011110011011",
    "1111100101011101",
    "1111110001010000",
    "1111111111111101",
    "1111110000011100",
    "1111100001111110",
    "1111010110010000",
    "1111001110101101",
    "1111001100100000",
    "1111010000010101",
    "1111011010001011",
    "1111101000111011",
    "1111111010100100",
    "1111110011100011",
    "1111100100001101",
    "1111011001011110",
    "1111010100100101",
    "1111010101110010",
    "1111011100101110",
    "1111101000111111",
    "1111111010001101",
    "1111110000010010",
    "1111011000001001",
    "1110111111110101",
    "1110101010100000",
    "1110011011000010",
    "1110010011010000",
    "1110010011010111",
    "1110011001111101",
    "1110100100100010",
    "1110110000001111",
    "1110111010100110",
    "1111000010000101",
    "1111000110010000",
    "1111000111101101",
    "1111000111111110",
    "1111001001001100",
    "1111001101110011",
    "1111010111101111",
    "1111100111110100",
    "1111111100111101",
    "1111101011101100",
    "1111010110001110",
    "1111000110100000",
    "1110111111000000",
    "1111000000000011",
    "1111000111101101",
    "1111010010101100",
    "1111011101101001",
    "1111100110001011",
    "1111101011110011",
    "1111110001011110",
    "1111111011111110",
    "1111110001000010",
    "1111010101011010",
    "1110110100111001",
    "1110010101110111",
    "1101111110110001",
    "1101110100001000",
    "1101110110110001",
    "1110000011101100",
    "1110010110110001",
    "1110101100100001",
    "1111000011010101",
    "1111011010111000",
    "1111110010100111",
    "1111110110111111",
    "1111100100011000",
    "1111011000100010",
    "1111010101111011",
    "1111011101100110",
    "1111101111000101",
    "1111111000000000",
    "1111011011110000",
    "1111000000100001",
    "1110101010000001",
    "1110011010101101",
    "1110010011101110",
    "1110010101011011",
    "1110011111111011",
    "1110110010110011",
    "1111001100111010",
    "1111101011110001",
    "1111110100010111",
    "1111011000000001",
    "1111000011000001",
    "1110110111110001",
    "1110110110010110",
    "1110111100111000",
    "1111001000101010",
    "1111010111101100",
    "1111101001101110",
    "1111111111101110",
    "1111100101011010",
    "1111000110011011",
    "1110100110001110",
    "1110001001011000",
    "1101110100101010",
    "1101101011001111",
    "1101101101100100",
    "1101111001111111",
    "1110001110001100",
    "1110101000011011",
    "1111000111111111",
    "1111101100010111",
    "1111101100001001",
    "1111000101000000",
    "1110100010100111",
    "1110001001011001",
    "1101111100000111",
    "1101111010111100",
    "1110000011011100",
    "1110010001110001",
    "1110100010010000",
    "1110110010011101",
    "1111000001100010",
    "1111001111101001",
    "1111011101001010",
    "1111101010000110",
    "1111110101110000",
    "1111111111001110",
    "1111111010000111",
    "1111110110010011",
    "1111110100100110",
    "1111110100000101",
    "1111110100001000",
    "1111110100101001",
    "1111110101111111",
    "1111111000010011",
    "1111111010111010",
    "1111111100001101",
    "1111111001111000",
    "1111110001101111",
    "1111100010101110",
    "1111001101101000",
    "1110110100111110",
    "1110011100100110",
    "1110001000100111",
    "1101111100000111",
    "1101111000100111",
    "1101111101100011",
    "1110001000111111",
    "1110011000010110",
    "1110101001000111",
    "1110111001011001",
    "1111001000110111",
    "1111011001000100",
    "1111101100010111",
    "1111111100000000",
    "1111100001001100",
    "1111000110101111",
    "1110110001111000",
    "1110100111110010",
    "1110101100001010",
    "1110111111001111",
    "1111011101010110",
    "1111111111100101",
    "1111011110010111",
    "1111000100001000",
    "1110110011010101",
    "1110101011110010",
    "1110101011001110",
    "1110101110011011",
    "1110110010110100",
    "1110110110111110",
    "1110111010100010",
    "1110111110000101",
    "1111000010010111",
    "1111001000000001",
    "1111001111101110",
    "1111011010001100",
    "1111101000001000",
    "1111111001101100",
    "1111110001110000",
    "1111011011110010",
    "1111000110001101",
    "1110110011000000",
    "1110100011110100",
    "1110011001011001",
    "1110010011100010",
    "1110010001000101",
    "1110010000110110",
    "1110010011000001",
    "1110011001100011",
    "1110100110100000",
    "1110111010011110",
    "1111010011011100",
    "1111101100101011",
    "1111111111010001",
    "1111110100111101",
    "1111110101111010",
    "1111111111111100",
    "1111110001000100",
    "1111100001111110",
    "1111010101011101",
    "1111001011101111",
    "1111000011011111",
    "1110111011011011",
    "1110110011010011",
    "1110101100100000",
    "1110101001011101",
    "1110101100101011",
    "1110110111110111",
    "1111001011010100",
    "1111100101101010",
    "1111111011110011",
    "1111011100011100",
    "1110111111101000",
    "1110101000011010",
    "1110011001011001",
    "1110010100010011",
    "1110011001010110",
    "1110100111011000",
    "1110111100100000",
    "1111010110100101",
    "1111110011101111",
    "1111101101100100",
    "1111001111000101",
    "1110110010101100",
    "1110011010100000",
    "1110001000100011",
    "1101111110011011",
    "1101111100101010",
    "1110000010101011",
    "1110001110111111",
    "1110011111010100",
    "1110110001011001",
    "1111000011001000",
    "1111010011000110",
    "1111100000011111",
    "1111101011000111",
    "1111110011000000",
    "1111111000011000",
    "1111111011010011",
    "1111111011111011",
    "1111111010101100",
    "1111111000010011",
    "1111110101111001",
    "1111110100101001",
    "1111110101100100",
    "1111111001001101",
    "1111111111100010",
    "1111110111111100",
    "1111101110010000",
    "1111100100011000",
    "1111011011010011",
    "1111010011100110",
    "1111001101100100",
    "1111001001010101",
    "1111000110110001",
    "1111000101101111",
    "1111000110001110",
    "1111001000011011",
    "1111001100110111",
    "1111010100110110",
    "1111100010001010",
    "1111110101110001",
    "1111110000101011",
    "1111010011011101",
    "1110110110010000",
    "1110011101000010",
    "1110001011000100",
    "1110000010000011",
    "1110000001100110",
    "1110000111110010",
    "1110010010001011",
    "1110011110010010",
    "1110101010001011",
    "1110110100100010",
    "1110111100101101",
    "1111000010101100",
    "1111000111111001",
    "1111001110101101",
    "1111011001100000",
    "1111101001001110",
    "1111111100100100",
    "1111101111101101",
    "1111100000000000",
    "1111011000010110",
    "1111011010111111",
    "1111100111010001",
    "1111111001110001",
    "1111110010011111",
    "1111100010011111",
    "1111011001111001",
    "1111011010100011",
    "1111100100010101",
    "1111110101000111",
    "1111110110100000",
    "1111100010011100",
    "1111010001111001",
    "1111000110110111",
    "1111000001111000",
    "1111000010010000",
    "1111000110100101",
    "1111001101011110",
    "1111010110000011",
    "1111100000001000",
    "1111101011111000",
    "1111111001001111",
    "1111111000011000",
    "1111101010001100",
    "1111011101011011",
    "1111010011000011",
    "1111001011011110",
    "1111000110010011",
    "1111000010100110",
    "1110111111010001",
    "1110111011100110",
    "1110110111110010",
    "1110110100110111",
    "1110110100001011",
    "1110110110110010",
    "1110111101000101",
    "1111000110100010",
    "1111010001100100",
    "1111011100011100",
    "1111100110101001",
    "1111110001010111",
    "1111111110010101",
    "1111110001100010",
    "1111011111101000",
    "1111001111000111",
    "1111000011111100",
    "1111000001001111",
    "1111000111110010",
    "1111010101100111",
    "1111100110111101",
    "1111111000001000",
    "1111111001000011",
    "1111101100110111",
    "1111100010001011",
    "1111011000000110",
    "1111001110101000",
    "1111000111001011",
    "1111000011111110",
    "1111000110110111",
    "1111010000101011",
    "1111100001000000",
    "1111110110011010",
    "1111110001000100",
    "1111010111100011",
    "1110111110111101",
    "1110101001001011",
    "1110011000001000",
    "1110001101010111",
    "1110001001100101",
    "1110001100001100",
    "1110010011011100",
    "1110011100110101",
    "1110100110000000",
    "1110101101001110",
    "1110110001100110",
    "1110110011001010",
    "1110110010011001",
    "1110110000000010",
    "1110101100110000",
    "1110101001000111",
    "1110100101110100",
    "1110100011101110",
    "1110100100000001",
    "1110101000000110",
    "1110110001001100",
    "1110111111110011",
    "1111010011010010",
    "1111101001110111",
    "1111111110110101",
    "1111101001010000",
    "1111010110111111",
    "1111001000101101",
    "1110111110000111",
    "1110110110100010",
    "1110110001010101",
    "1110101110001111",
    "1110101101100000",
    "1110101111110000",
    "1110110101101010",
    "1110111111011001",
    "1111001100100011",
    "1111011100001001",
    "1111101100110100",
    "1111111101000111",
    "1111110100010111",
    "1111101000101010",
    "1111100000000111",
    "1111011010100010",
    "1111010111011000",
    "1111010101111001",
    "1111010101010000",
    "1111010100110110",
    "1111010100000110",
    "1111010010110110",
    "1111010001000111",
    "1111001111010010",
    "1111001110001010",
    "1111001110101101",
    "1111010001110110",
    "1111010111111111",
    "1111100000110011",
    "1111101010111100",
    "1111110100100001",
    "1111111011101000",
    "1111111110110101",
    "1111111101110000",
    "1111111001001100",
    "1111110010111100",
    "1111101101001010",
    "1111101010000000",
    "1111101011001000",
    "1111110001100100",
    "1111111101011111",
    "1111110001111010",
    "1111011110011111",
    "1111001010101111",
    "1110111001001011",
    "1110101100000001",
    "1110100100100100",
    "1110100011000101",
    "1110100110110010",
    "1110101110001111",
    "1110110111110111",
    "1111000010100111",
    "1111001110010100",
    "1111011011010100",
    "1111101010000110",
    "1111111010011001",
    "1111110101001010",
    "1111100111000000",
    "1111011101110011",
    "1111011011101000",
    "1111100000111101",
    "1111101100010000",
    "1111111010101001",
    "1111110111010000",
    "1111101100001101",
    "1111100101011000",
    "1111100010011101",
    "1111100001110000",
    "1111100001000010",
    "1111011110010110",
    "1111011000100011",
    "1111001111101001",
    "1111000100101001",
    "1110111001000110",
    "1110101110110101",
    "1110100111100111",
    "1110100100101100",
    "1110100110100111",
    "1110101100111010",
    "1110110110010011",
    "1111000001000111",
    "1111001011101000",
    "1111010101000000",
    "1111011110001100",
    "1111101001100011",
    "1111111001100101",
    "1111110000110110",
    "1111010111100000",
    "1110111110010001",
    "1110101001101111",
    "1110011101011110",
    "1110011010101111",
    "1110011111110000",
    "1110101000111111",
    "1110110011000001",
    "1110111011111111",
    "1111000100011100",
    "1111001110001001",
    "1111011010110111",
    "1111101010111110",
    "1111111100110111",
    "1111110010011101",
    "1111100110011011",
    "1111100001001111",
    "1111100011010000",
    "1111101010110000",
    "1111110101000001",
    "1111111111010110",
    "1111110111111111",
    "1111110001110010",
    "1111101110000001",
    "1111101100100000",
    "1111101101000001",
    "1111101111010101",
    "1111110011000001",
    "1111110111011010",
    "1111111011100111",
    "1111111110101001",
    "1111111111101100",
    "1111111110011000",
    "1111111010111000",
    "1111110101101111",
    "1111101111100000",
    "1111101000100110",
    "1111100001010010",
    "1111011001100101",
    "1111010001010101",
    "1111001000101000",
    "1110111111100110",
    "1110110110100111",
    "1110101110000111",
    "1110100110100010",
    "1110100000010111",
    "1110011100010001",
    "1110011011000010",
    "1110011101011011",
    "1110100011111011",
    "1110101110101011",
    "1110111101010010",
    "1111001110111010",
    "1111100010001010",
    "1111110101011101",
    "1111111000110000",
    "1111101001111100",
    "1111011111000000",
    "1111011000011011",
    "1111010110010010",
    "1111011000001001",
    "1111011101011100",
    "1111100101011010",
    "1111101111011011",
    "1111111010111010",
    "1111111000101111",
    "1111101100011000",
    "1111100000111110",
    "1111010111100011",
    "1111010001001000",
    "1111001110101000",
    "1111010000101011",
    "1111010111100010",
    "1111100010110011",
    "1111110001001001",
    "1111111111100101",
    "1111110010001100",
    "1111101001011100",
    "1111100111100101",
    "1111101101111011",
    "1111111100011101",
    "1111101110010110",
    "1111010101100111",
    "1110111101001100",
    "1110101000111111",
    "1110011011111010",
    "1110010111011011",
    "1110011011010001",
    "1110100101111011",
    "1110110101100111",
    "1111001001000100",
    "1111011111101100",
    "1111111001001001",
    "1111101011101001",
    "1111010000111110",
    "1110111001111100",
    "1110101001101000",
    "1110100010001011",
    "1110100100000011",
    "1110101101111101",
    "1110111101010010",
    "1111001111001010",
    "1111100001000011",
    "1111110001010010",
    "1111111110111011",
    "1111110110011100",
    "1111101111000101",
    "1111101010111010",
    "1111101001011000",
    "1111101001011100",
    "1111101001101111",
    "1111101001001110",
    "1111100111101011",
    "1111100101110110",
    "1111100101001110",
    "1111100111010111",
    "1111101101001100",
    "1111110110110001",
    "1111111100101000",
    "1111101110011011",
    "1111100000000111",
    "1111010011001010",
    "1111001000111010",
    "1111000010011100",
    "1111000000010100",
    "1111000010110011",
    "1111001001110000",
    "1111010100110011",
    "1111100011010101",
    "1111110100011111",
    "1111111001000111",
    "1111100111100100",
    "1111011001000110",
    "1111001111100011",
    "1111001011110011",
    "1111001101100011",
    "1111010011010101",
    "1111011011000110",
    "1111100010111011",
    "1111101001111000",
    "1111110000001000",
    "1111110110110001",
    "1111111111001000",
    "1111110101111110",
    "1111101000111110",
    "1111011011101000",
    "1111010000101011",
    "1111001010110101",
    "1111001100010011",
    "1111010101111011",
    "1111100111000100",
    "1111111101011011",
    "1111101010011111",
    "1111010100101100",
    "1111000100100000",
    "1110111100000010",
    "1110111011110011",
    "1111000010111001",
    "1111001111101001",
    "1111100000001111",
    "1111110011011001",
    "1111110111110100",
    "1111100010100100",
    "1111001110010111",
    "1110111101010110",
    "1110110001100001",
    "1110101100100110",
    "1110101111011001",
    "1110111001110010",
    "1111001010100101",
    "1111011111110101",
    "1111110110110111",
    "1111110010111100",
    "1111011111110001",
    "1111010000111011",
    "1111000110101101",
    "1111000000110011",
    "1110111110001111",
    "1110111110000010",
    "1110111111011010",
    "1111000010001000",
    "1111000110011000",
    "1111001100011001",
    "1111010100010101",
    "1111011101111000",
    "1111101000010100",
    "1111110010100001",
    "1111111011001011",
    "1111111110110011",
    "1111111100001100",
    "1111111100111110",
    "1111111111010100",
    "1111111001110010",
    "1111110011101001",
    "1111101110001111",
    "1111101010101010",
    "1111101001101011",
    "1111101011100111",
    "1111110000011111",
    "1111111000001001",
    "1111111101100100",
    "1111110000111010",
    "1111100001111110",
    "1111010000111011",
    "1110111110001111",
    "1110101010111111",
    "1110011000110010",
    "1110001001101011",
    "1101111111100100",
    "1101111011100110",
    "1101111101110010",
    "1110000100110001",
    "1110001110010111",
    "1110011000001110",
    "1110100000100111",
    "1110100111110001",
    "1110101111100001",
    "1110111001111001",
    "1111000111011111",
    "1111010110010101",
    "1111100010010100",
    "1111100110100010",
    "1111011111010010",
    "1111001011111010",
    "1110101111101001",
    "1110010000101001",
    "1101110101101111",
    "1101100100000101",
    "1101011101101001",
    "1101100001011100",
    "1101101101010100",
    "1101111111111111",
    "1110011000111111",
    "1110110111110101",
    "1111011010100011",
    "1111111101011010",
    "1111100100001011",
    "1111001110110000",
    "1111000100110111",
    "1111000101101110",
    "1111001101011001",
    "1111010110111110",
    "1111011110010010",
    "1111100001100100",
    "1111100001010101",
    "1111011111110000",
    "1111011111101001",
    "1111100011010101",
    "1111101011110111",
    "1111111000111001",
    "1111110110101110",
    "1111100100110001",
    "1111010010110110",
    "1111000010100001",
    "1110110101001011",
    "1110101100000010",
    "1110100111111001",
    "1110101000101000",
    "1110101101000101",
    "1110110011011100",
    "1110111001101111",
    "1110111110011001",
    "1111000000101001",
    "1111000000100100",
    "1110111111001100",
    "1110111110010100",
    "1110111111111011",
    "1111000101001101",
    "1111001110000010",
    "1111011001000001",
    "1111100011110100",
    "1111101011110011",
    "1111101110110111",
    "1111101100001011",
    "1111100100010011",
    "1111011000111010",
    "1111001100010111",
    "1111000001010100",
    "1110111010010100",
    "1110111001010001",
    "1110111111001100",
    "1111001100010110",
    "1111100000100110",
    "1111111011001111",
    "1111100101011010",
    "1111000100010101",
    "1110100101010111",
    "1110001100010110",
    "1101111100000101",
    "1101110101100111",
    "1101111000000011",
    "1110000001001010",
    "1110001110100011",
    "1110011110101001",
    "1110110000111011",
    "1111000101001110",
    "1111011010111111",
    "1111110000101011",
    "1111111011111101",
    "1111101101011011",
    "1111100101011101",
    "1111100100010010",
    "1111101000101000",
    "1111110000001001",
    "1111111000011110",
    "1111111111111100",
    "1111111001101011",
    "1111110100010110",
    "1111101111100011",
    "1111101011011010",
    "1111101000101110",
    "1111101000101000",
    "1111101100000101",
    "1111110011010110",
    "1111111101110100",
    "1111110101101111",
    "1111101000111111",
    "1111011101001111",
    "1111010011011010",
    "1111001100000010",
    "1111000111100000",
    "1111000110010101",
    "1111001001110100",
    "1111010011101001",
    "1111100101000101",
    "1111111101101011",
    "1111100100111110",
    "1111000111000011",
    "1110101101010100",
    "1110011011101101",
    "1110010100001000",
    "1110010110001000",
    "1110011111010110",
    "1110101100110101",
    "1110111100001111",
    "1111001100010110",
    "1111011100110101",
    "1111101101100100",
    "1111111101111110",
    "1111110011010000",
    "1111101000000101",
    "1111100010001011",
    "1111100010011111",
    "1111101001000010",
    "1111110101001011",
    "1111111001101111",
    "1111100100000101",
    "1111001010001001",
    "1110101101000111",
    "1110001111001111",
    "1101110011111001",
    "1101011110100110",
    "1101010010001111",
    "1101010000010010",
    "1101011000110101",
    "1101101010111111",
    "1110000101010011",
    "1110100101101001",
    "1111001001000010",
    "1111101011101111",
    "1111110110011011",
    "1111100001010111",
    "1111010111101101",
    "1111011010011000",
    "1111101000101010",
    "1111111111100101",
    "1111100001110011",
    "1111000010000101",
    "1110100100100111",
    "1110001101000000",
    "1101111101101110",
    "1101110111111001",
    "1101111011011000",
    "1110000111000100",
    "1110011001010101",
    "1110110000001000",
    "1111001001001100",
    "1111100010000010",
    "1111111000001001",
    "1111110110100010",
    "1111101011011111",
    "1111100111001000",
    "1111101000111111",
    "1111101111100010",
    "1111111000110011",
    "1111111101010000",
    "1111110100011110",
    "1111101101110111",
    "1111101001101001",
    "1111100111001011",
    "1111100101100000",
    "1111100011111000",
    "1111100001111011",
    "1111011111110011",
    "1111011101111000",
    "1111011100100000",
    "1111011011100101",
    "1111011010101000",
    "1111011001001110",
    "1111010111010000",
    "1111010101000001",
    "1111010011100010",
    "1111010011110011",
    "1111010110011101",
    "1111011011101000",
    "1111100010110110",
    "1111101011101000",
    "1111110101111100",
    "1111111101110100",
    "1111101111010110",
    "1111011110111101",
    "1111001101111010",
    "1110111110001101",
    "1110110010000000",
    "1110101010110000",
    "1110101000111110",
    "1110101100000100",
    "1110110011001011",
    "1110111101110111",
    "1111001100001100",
    "1111011110011110",
    "1111110100001101",
    "1111110100001011",
    "1111011101100001",
    "1111001011000111",
    "1110111111110000",
    "1110111100110000",
    "1111000001011010",
    "1111001011001100",
    "1111010110110001",
    "1111100000111011",
    "1111100111011011",
    "1111101001011011",
    "1111100111001011",
    "1111100001101100",
    "1111011010010011",
    "1111010010010010",
    "1111001010101000",
    "1111000100000110",
    "1110111111000111",
    "1110111100001001",
    "1110111011101111",
    "1110111110011011",
    "1111000100110001",
    "1111001111000000",
    "1111011100111000",
    "1111101101100000",
    "1111111111011001",
    "1111101111001111",
    "1111100000010010",
    "1111010101010000",
    "1111001111010100",
    "1111001110111111",
    "1111010100001011",
    "1111011110000111",
    "1111101011010011",
    "1111111001111111",
    "1111110111011101",
    "1111101010011011",
    "1111011111101000",
    "1111010111010110",
    "1111010001110000",
    "1111001110110110",
    "1111001110111000",
    "1111010010000010",
    "1111011000010011",
    "1111100001010100",
    "1111101100010100",
    "1111111000011010",
    "1111111011001110",
    "1111101111001011",
    "1111100011100010",
    "1111011000010011",
    "1111001101010110",
    "1111000010111001",
    "1110111001100101",
    "1110110010010111",
    "1110101110001001",
    "1110101101011001",
    "1110110000000000",
    "1110110101010000",
    "1110111011111101",
    "1111000010110100",
    "1111001000011010",
    "1111001011100000",
    "1111001011001010",
    "1111000110110110",
    "1110111110011110",
    "1110110010101100",
    "1110100100110110",
    "1110010110111100",
    "1110001011001010",
    "1110000011100111",
    "1110000001111011",
    "1110000111001001",
    "1110010011111001",
    "1110101000011101",
    "1111000100011000",
    "1111100110000001",
    "1111110101110011",
    "1111010011100111",
    "1110110111110101",
    "1110100101110100",
    "1110011110110001",
    "1110100001011100",
    "1110101010110101",
    "1110110111011011",
    "1111000100011100",
    "1111010000011111",
    "1111011011100101",
    "1111100110001101",
    "1111110000100111",
    "1111111010011010",
    "1111111101010001",
    "1111110111011010",
    "1111110100010000",
    "1111110011000100",
    "1111110001111110",
    "1111101110011101",
    "1111100101111100",
    "1111010111000001",
    "1111000010001011",
    "1110101001111001",
    "1110010001110100",
    "1101111101111000",
    "1101110001001000",
    "1101101100110111",
    "1101110000011001",
    "1101111001010110",
    "1110000100110111",
    "1110010001010100",
    "1110011111110011",
    "1110110010111011",
    "1111001100110011",
    "1111101101000111",
    "1111101111101000",
    "1111001111001000",
    "1110110111001110",
    "1110101011110010",
    "1110101101000101",
    "1110110111111110",
    "1111000111111010",
    "1111011001000100",
    "1111101001111100",
    "1111111011010000",
    "1111110001110101",
    "1111011101000111",
    "1111001000000011",
    "1110110101101100",
    "1110101001101000",
    "1110100110011010",
    "1110101100101011",
    "1110111011000010",
    "1111001110011110",
    "1111100011100111",
    "1111110111100001",
    "1111111000000010",
    "1111101100111100",
    "1111101000101001",
    "1111101100001001",
    "1111110111010101",
    "1111110111001111",
    "1111100010010111",
    "1111001101011110",
    "1110111011111010",
    "1110110000001010",
    "1110101011101010",
    "1110101110101011",
    "1110111001000001",
    "1111001010000111",
    "1111100001001100",
    "1111111100101101",
    "1111100101101100",
    "1111001001010101",
    "1110110001010101",
    "1110100000001101",
    "1110010110111110",
    "1110010100111100",
    "1110011000010011",
    "1110011110111010",
    "1110100111011011",
    "1110110001110000",
    "1110111110100110",
    "1111001110111101",
    "1111100011000000",
    "1111111001111000",
    "1111101110001010",
    "1111010111010110",
    "1111000011101001",
    "1110110100010010",
    "1110101001101111",
    "1110100011101001",
    "1110100001010100",
    "1110100001111110",
    "1110100100111011",
    "1110101001001011",
    "1110101101101110",
    "1110110001101100",
    "1110110100100100",
    "1110110110010011",
    "1110110111100000",
    "1110111001000001",
    "1110111011101111",
    "1111000000001100",
    "1111000110010011",
    "1111001101011110",
    "1111010100101111",
    "1111011011010011",
    "1111100000101110",
    "1111100101001110",
    "1111101001011111",
    "1111101110011100",
    "1111110101001010",
    "1111111110101011",
    "1111110100000111",
    "1111100011000001",
    "1111001110110110",
    "1110111001110000",
    "1110100110110110",
    "1110011001000110",
    "1110010010100111",
    "1110010011110001",
    "1110011011010110",
    "1110100110111001",
    "1110110011111110",
    "1111000001000000",
    "1111001101101011",
    "1111011010011000",
    "1111100111010010",
    "1111110011100110",
    "1111111101010110",
    "1111111101111111",
    "1111111111010101",
    "1111110100110100",
    "1111100011110100",
    "1111001111011001",
    "1110111011010110",
    "1110101011000010",
    "1110100000010100",
    "1110011011010011",
    "1110011011000001",
    "1110011101110111",
    "1110100010010111",
    "1110100111010000",
    "1110101011100110",
    "1110101110101110",
    "1110110000010101",
    "1110110000011111",
    "1110101111110110",
    "1110101111101001",
    "1110110001111000",
    "1110111000110100",
    "1111000110011000",
    "1111011011010110",
    "1111110110100010",
    "1111101011001100",
    "1111001110001010",
    "1110110110010101",
    "1110100110010011",
    "1110011110100011",
    "1110011101100001",
    "1110100000011110",
    "1110100100100010",
    "1110101000000110",
    "1110101011100101",
    "1110110001001000",
    "1110111011001001",
    "1111001010100101",
    "1111011110001111",
    "1111110010110110",
    "1111111011110010",
    "1111110001011100",
    "1111101111111010",
    "1111110110101000",
    "1111111100111000",
    "1111101101111110",
    "1111011111101100",
    "1111010100011000",
    "1111001101011001",
    "1111001011011000",
    "1111001110011110",
    "1111010110101100",
    "1111100100010010",
    "1111110111011111",
    "1111110000001110",
    "1111010100101100",
    "1110111000111111",
    "1110100001000011",
    "1110010000010101",
    "1110001000111100",
    "1110001010111000",
    "1110010100010111",
    "1110100010001111",
    "1110110001010100",
    "1110111111000010",
    "1111001010111111",
    "1111010111001101",
    "1111100110101001",
    "1111111011011011",
    "1111101010101100",
    "1111001110111000",
    "1110110101110100",
    "1110100100010010",
    "1110011101010111",
    "1110100000110101",
    "1110101011100011",
    "1110111001000111",
    "1111000101011111",
    "1111001110001111",
    "1111010010110001",
    "1111010100000001",
    "1111010011110110",
    "1111010011111100",
    "1111010101000011",
    "1111010110110001",
    "1111010111110111",
    "1111010111000110",
    "1111010011111000",
    "1111001110011111",
    "1111000111111100",
    "1111000001011100",
    "1110111100001111",
    "1110111001110000",
    "1110111011011110",
    "1111000010010010",
    "1111001101111011",
    "1111011100110111",
    "1111101100011010",
    "1111111001110000",
    "1111111101010000",
    "1111111001100010",
    "1111111010001010",
    "1111111100111111",
    "1111111111101101",
    "1111111111010011",
    "1111111111100010",
    "1111111101010001",
    "1111111011101100",
    "1111111100110111",
    "1111111101101110",
    "1111110100000111",
    "1111100111101101",
    "1111011011000001",
    "1111010000101011",
    "1111001010110101",
    "1111001010110000",
    "1111010000111000",
    "1111011100111111",
    "1111101110100100",
    "1111111010110110",
    "1111100000010101",
    "1111000011110001",
    "1110101000001001",
    "1110010000111110",
    "1110000001011001",
    "1101111011001001",
    "1101111110001111",
    "1110001001010101",
    "1110011010011110",
    "1110101111110110",
    "1111000111110010",
    "1111100000011111",
    "1111110111111111",
    "1111110100000011",
    "1111100101110111",
    "1111011110110000",
    "1111011110101110",
    "1111100100100100",
    "1111101110001011",
    "1111111001011101",
    "1111111011000001",
    "1111110000001001",
    "1111100110001110",
    "1111011101101000",
    "1111010110111110",
    "1111010010111110",
    "1111010010001101",
    "1111010100100000",
    "1111011000110111",
    "1111011101101101",
    "1111100001100100",
    "1111100011101110",
    "1111100100100101",
    "1111100101011000",
    "1111100111101111",
    "1111101100101011",
    "1111110100010111",
    "1111111101101110",
    "1111111001000010",
    "1111110010000110",
    "1111101111010001",
    "1111110001100010",
    "1111111001000101",
    "1111111010011101",
    "1111101001110001",
    "1111010101100100",
    "1110111111000111",
    "1110101000011011",
    "1110010100000011",
    "1110000100100100",
    "1101111011110101",
    "1101111010101000",
    "1110000000001101",
    "1110001010100101",
    "1110010111010101",
    "1110100100100111",
    "1110110010001101",
    "1111000001011100",
    "1111010100001110",
    "1111101011100111",
    "1111111001001100",
    "1111011101010110",
    "1111000101001000",
    "1110110100100101",
    "1110101110000100",
    "1110110001010100",
    "1110111011111101",
    "1111001010110101",
    "1111011011010100",
    "1111101100010100",
    "1111111101111010",
    "1111101111100001",
    "1111011100010110",
    "1111001001111010",
    "1110111010101000",
    "1110110001000011",
    "1110101110111010",
    "1110110100001000",
    "1110111110101101",
    "1111001011001110",
    "1111010110001000",
    "1111011100101101",
    "1111011101100110",
    "1111011000111001",
    "1111001111101100",
    "1111000011110011",
    "1110110111001001",
    "1110101011101010",
    "1110100010111000",
    "1110011101101101",
    "1110011100010011",
    "1110011101111111",
    "1110100001101100",
    "1110100110011011",
    "1110101100000101",
    "1110110011101111",
    "1110111111000101",
    "1111001111011110",
    "1111100101000110",
    "1111111110100101",
    "1111100110111100",
    "1111001111000010",
    "1110111100100001",
    "1110110000110110",
    "1110101011110000",
    "1110101011111111",
    "1110110000000111",
    "1110110111001000",
    "1111000000100011",
    "1111001011111111",
    "1111011000110000",
    "1111100101100100",
    "1111110000101100",
    "1111111000011111",
    "1111111100000001",
    "1111111011011001",
    "1111110111110101",
    "1111110011000111",
    "1111101110101101",
    "1111101011010100",
    "1111101000101000",
    "1111100101100100",
    "1111100000101110",
    "1111011001000111",
    "1111001110101110",
    "1111000010100100",
    "1110110110100000",
    "1110101100101000",
    "1110100110101101",
    "1110100110001110",
    "1110101100001111",
    "1110111001100011",
    "1111001110001100",
    "1111101000101110",
    "1111111001111111",
    "1111011110011011",
    "1111001000111110",
    "1110111100111111",
    "1110111011101011",
    "1111000100000001",
    "1111010011100010",
    "1111100111011110",
    "1111111101110001",
    "1111101010111110",
    "1111010100011010",
    "1111000000101001",
    "1110110010010111",
    "1110101100010111",
    "1110110000111001",
    "1111000000110001",
    "1111011010100011",
    "1111111010010001",
    "1111100101011000",
    "1111001001110000",
    "1110110110011010",
    "1110101100101000",
    "1110101011100000",
    "1110110000100011",
    "1110111000110000",
    "1111000001111000",
    "1111001010111111",
    "1111010100100010",
    "1111011111110001",
    "1111101101101110",
    "1111111110011110",
    "1111101111000011",
    "1111011101000010",
    "1111001101111000",
    "1111000011011000",
    "1110111110000111",
    "1110111101001110",
    "1110111110111011",
    "1111000001101011",
    "1111000100011111",
    "1111000111010011",
    "1111001010011000",
    "1111001110001100",
    "1111010011001000",
    "1111011001101010",
    "1111100001111001",
    "1111101011101110",
    "1111110110011110",
    "1111111110110010",
    "1111110101010010",
    "1111101110000000",
    "1111101001100001",
    "1111100111110100",
    "1111101000010010",
    "1111101001111101",
    "1111101011111100",
    "1111101101101010",
    "1111101110111110",
    "1111110000000010",
    "1111110001000000",
    "1111110001111001",
    "1111110010110011",
    "1111110011111010",
    "1111110101101100",
    "1111111000110000",
    "1111111101100110",
    "1111111011110011",
    "1111110100011000",
    "1111101101011111",
    "1111101000100101",
    "1111100110100011",
    "1111100111010001",
    "1111101001110000",
    "1111101100010101",
    "1111101101010011",
    "1111101011011110",
    "1111100110100101",
    "1111011111010001",
    "1111010110111110",
    "1111001111001111",
    "1111001001011000",
    "1111000110001001",
    "1111000101100100",
    "1111000111001000",
    "1111001001111100",
    "1111001101000100",
    "1111001111100011",
    "1111010000110000",
    "1111010000001100",
    "1111001101101011",
    "1111001001010110",
    "1111000011100001",
    "1110111100101011",
    "1110110101010011",
    "1110101101111000",
    "1110100110110111",
    "1110100000101011",
    "1110011011100011",
    "1110010111100011",
    "1110010100100101",
    "1110010010010111",
    "1110010000101011",
    "1110001111010111",
    "1110001110101001",
    "1110001111000100",
    "1110010001001000",
    "1110010101010011",
    "1110011011011101",
    "1110100010110001",
    "1110101010000001",
    "1110101111110110",
    "1110110011010010",
    "1110110100001000",
    "1110110011000000",
    "1110110001001000",
    "1110101111111011",
    "1110110000100100",
    "1110110011110011",
    "1110111001100101",
    "1111000001010100",
    "1111001001111100",
    "1111010010001010",
    "1111011000110010",
    "1111011100111101",
    "1111011110010111",
    "1111011101010010",
    "1111011010100000",
    "1111010111001101",
    "1111010100101111",
    "1111010100011101",
    "1111010111100101",
    "1111011111000010",
    "1111101011010101",
    "1111111100001101",
    "1111101111101010",
    "1111011010110111",
    "1111001000011101",
    "1110111011010110",
    "1110110101011111",
    "1110110111100000",
    "1111000000111000",
    "1111010000010010",
    "1111100011111100",
    "1111111001110010",
    "1111110000110001",
    "1111011110100100",
    "1111010010011001",
    "1111001110011100",
    "1111010100001010",
    "1111100011100111",
    "1111111011011110",
    "1111100111000101",
    "1111000111111010",
    "1110101010110111",
    "1110010011001010",
    "1110000010101111",
    "1101111010011000",
    "1101111001100101",
    "1101111111010001",
    "1110001010000111",
    "1110011000110101",
    "1110101001111010",
    "1110111011100000",
    "1111001011100110",
    "1111011000010110",
    "1111100000100011",
    "1111100100000000",
    "1111100011101110",
    "1111100001101011",
    "1111100000011110",
    "1111100010100001",
    "1111101001001111",
    "1111110100010100",
    "1111111110001110",
    "1111110001001111",
    "1111100111011000",
    "1111100010001111",
    "1111100001111101",
    "1111100101011011",
    "1111101010100111",
    "1111101111011001",
    "1111110010001000",
    "1111110010001001",
    "1111110000000011",
    "1111101101111001",
    "1111101110110001",
    "1111110101100011",
    "1111111100011001",
    "1111101000000010",
    "1111010000011010",
    "1110111001110101",
    "1110101000010110",
    "1110011110011110",
    "1110011100011100",
    "1110100000100110",
    "1110101000011101",
    "1110110001110011",
    "1110111011011110",
    "1111000101010101",
    "1111001111101000",
    "1111011010010100",
    "1111100100011101",
    "1111101100011101",
    "1111110000100010",
    "1111101111101000",
    "1111101001111111",
    "1111100001001101",
    "1111010111110010",
    "1111010000010100",
    "1111001100110011",
    "1111001110010001",
    "1111010100100100",
    "1111011110100100",
    "1111101010011111",
    "1111110110010100",
    "1111111111101000",
    "1111111000100001",
    "1111110100101010",
    "1111110011110000",
    "1111110100111111",
    "1111110111011000",
    "1111111010001010",
    "1111111101000001",
    "1111111111110000",
    "1111111011100111",
    "1111110101110101",
    "1111101110000001",
    "1111100100011000",
    "1111011001101011",
    "1111001111001111",
    "1111000110011101",
    "1111000000100111",
    "1110111110100110",
    "1111000000110101",
    "1111000111011000",
    "1111010001111101",
    "1111011111110001",
    "1111101111101000",
    "1111111111101110",
    "1111110001111010",
    "1111100111010010",
    "1111100001110011",
    "1111100001111001",
    "1111100111000001",
    "1111101111100111",
    "1111111001110101",
    "1111111011111001",
    "1111110010100000",
    "1111101010000101",
    "1111100010001011",
    "1111011010010011",
    "1111010010001010",
    "1111001001111001",
    "1111000010000000",
    "1110111011001111",
    "1110110110010110",
    "1110110100000001",
    "1110110100111011",
    "1110111001100111",
    "1111000010010010",
    "1111001110100100",
    "1111011101000101",
    "1111101011100001",
    "1111110111000111",
    "1111111101010101",
    "1111111100100101",
    "1111110100100111",
    "1111100110100110",
    "1111010101000101",
    "1111000011011101",
    "1110110101011101",
    "1110101110011111",
    "1110110001000111",
    "1110111110011011",
    "1111010101100111",
    "1111110011110010",
    "1111101011011010",
    "1111001100111000",
    "1110110100110001",
    "1110100101100100",
    "1110011111100100",
    "1110100001001111",
    "1110100111110010",
    "1110110000110101",
    "1110111011100101",
    "1111001001011001",
    "1111011100010110",
    "1111110101011001",
    "1111101100111010",
    "1111001110101000",
    "1110110101000011",
    "1110100100111110",
    "1110100000110001",
    "1110100111001001",
    "1110110011111000",
    "1111000001011111",
    "1111001011001110",
    "1111001110100011",
    "1111001011011101",
    "1111000011110011",
    "1110111010100101",
    "1110110010100111",
    "1110101101101011",
    "1110101100010110",
    "1110101110011110",
    "1110110011111000",
    "1110111100110101",
    "1111001001111001",
    "1111011011000100",
    "1111101111001101",
    "1111111011110100",
    "1111101001000000",
    "1111011011001110",
    "1111010100111001",
    "1111010111000001",
    "1111100000101110",
    "1111101111101010",
    "1111111111011001",
    "1111101111101011",
    "1111100011011100",
    "1111011011101111",
    "1111011000010110",
    "1111011000010110",
    "1111011010101011",
    "1111011111000000",
    "1111100101110010",
    "1111101111111111",
    "1111111110001100",
    "1111101111111111",
    "1111011100011001",
    "1111001001110010",
    "1110111011000010",
    "1110110010011100",
    "1110110000101100",
    "1110110101000101",
    "1110111110001101",
    "1111001011000111",
    "1111011011101111",
    "1111110000001010",
    "1111111000010001",
    "1111011111111011",
    "1111001010100010",
    "1110111100010001",
    "1110111000011110",
    "1111000000101011",
    "1111010100001101",
    "1111110000011001",
    "1111101110110001",
    "1111001101101101",
    "1110110000000111",
    "1110011000110000",
    "1110001001000100",
    "1110000001010100",
    "1110000000111000",
    "1110000110101100",
    "1110010001110000",
    "1110100001011111",
    "1110110101011011",
    "1111001100111111",
    "1111100110111011",
    "1111111110100110",
    "1111100110000011",
    "1111010001111000",
    "1111000100001000",
    "1110111101101011",
    "1110111110001100",
    "1111000100001101",
    "1111001110000100",
    "1111011010011000",
    "1111101000010010",
    "1111110111000101",
    "1111111001111110",
    "1111101100010100",
    "1111100001100111",
    "1111011011101000",
    "1111011011100011",
    "1111100001100100",
    "1111101100101000",
    "1111111010100110",
    "1111110111001000",
    "1111101011010111",
    "1111100100001010",
    "1111100010101011",
    "1111100111000011",
    "1111110000100010",
    "1111111101110111",
    "1111110010001101",
    "1111100000101001",
    "1111001101110011",
    "1110111001110100",
    "1110100101010000",
    "1110010001010000",
    "1101111111101000",
    "1101110010011100",
    "1101101011101010",
    "1101101100011011",
    "1101110100111011",
    "1110000101000000",
    "1110011100100001",
    "1110111011001001",
    "1111011111100001",
    "1111111001011111",
    "1111010100100101",
    "1110110110101010",
    "1110100011101001",
    "1110011101001100",
    "1110100010001011",
    "1110101111001000",
    "1111000000000111",
    "1111010010100001",
    "1111100101101110",
    "1111111010010010",
    "1111101111011000",
    "1111011000011110",
    "1111000100000101",
    "1110110110100101",
    "1110110100100100",
    "1111000000010111",
    "1111011000110000",
    "1111111000111000",
    "1111100110001101",
    "1111001011001110",
    "1110111010100010",
    "1110110101011101",
    "1110111010011000",
    "1111000101110111",
    "1111010100101001",
    "1111100100011000",
    "1111110100010011",
    "1111111011011010",
    "1111101010101001",
    "1111011001110101",
    "1111001010001001",
    "1110111100111100",
    "1110110011010011",
    "1110101101011001",
    "1110101010101000",
    "1110101001110010",
    "1110101001110000",
    "1110101001111001",
    "1110101010001110",
    "1110101011001010",
    "1110101101000010",
    "1110101111110011",
    "1110110011010101",
    "1110111000001110",
    "1111000000000111",
    "1111001100101000",
    "1111011110100001",
    "1111110100011010",
    "1111110101000010",
    "1111100010011100",
    "1111010111111010",
    "1111010111100011",
    "1111100000100111",
    "1111110000000001",
    "1111111101111001",
    "1111101011111011",
    "1111011010101010",
    "1111001001010101",
    "1110110111010000",
    "1110100100101001",
    "1110010011010010",
    "1110000101110111",
    "1101111111000100",
    "1110000000001010",
    "1110001000011011",
    "1110010101010010",
    "1110100011101110",
    "1110110001111101",
    "1111000000010001",
    "1111010000011111",
    "1111100100011000",
    "1111111011111101",
    "1111101010110100",
    "1111010100000001",
    "1111000100000101",
    "1110111110000000",
    "1111000010011100",
    "1111001111000010",
    "1111011111110000",
    "1111110000000001",
    "1111111100001011",
    "1111111110000001",
    "1111111111010000",
    "1111111001001101",
    "1111101101001010",
    "1111011110100110",
    "1111001111011111",
    "1111000001100001",
    "1110110110000011",
    "1110101110000100",
    "1110101001110101",
    "1110101001000100",
    "1110101011000100",
    "1110101111101001",
    "1110110111101000",
    "1111000100100100",
    "1111010111011111",
    "1111110000000100",
    "1111110100000010",
    "1111011000101010",
    "1111000001110001",
    "1110110010011100",
    "1110101011101000",
    "1110101100101101",
    "1110110100010011",
    "1111000001011111",
    "1111010100000101",
    "1111101011111101",
    "1111110111111101",
    "1111011010010001",
    "1110111110100011",
    "1110101000101010",
    "1110011011100000",
    "1110011000001001",
    "1110011101101101",
    "1110101001101101",
    "1110111001010001",
    "1111001010001011",
    "1111011011001111",
    "1111101100010100",
    "1111111101011001",
    "1111110001111100",
    "1111100010110100",
    "1111010110100101",
    "1111001110100100",
    "1111001011100001",
    "1111001101011001",
    "1111010011100001",
    "1111011101000000",
    "1111101001010101",
    "1111111000011001",
    "1111110110001001",
    "1111100011100110",
    "1111010010000010",
    "1111000011111110",
    "1110111011101010",
    "1110111010011011",
    "1111000000100100",
    "1111001101010111",
    "1111011111100110",
    "1111110101111010",
    "1111110001001110",
    "1111011000001110",
    "1111000010001010",
    "1110110010100111",
    "1110101100101010",
    "1110110010000000",
    "1111000010100110",
    "1111011100110111",
    "1111111101110101",
    "1111011110001101",
    "1110111011100101",
    "1110011101111101",
    "1110001000001001",
    "1101111011100001",
    "1101111000001011",
    "1101111100111000",
    "1110000111110001",
    "1110010110110010",
    "1110101000100111",
    "1110111100101010",
    "1111010010101011",
    "1111101010000100",
    "1111111110010101",
    "1111101000010100",
    "1111010101100111",
    "1111000111011101",
    "1110111110001001",
    "1110111000110100",
    "1110110101111011",
    "1110110100000000",
    "1110110010010101",
    "1110110001001100",
    "1110110001001111",
    "1110110011000000",
    "1110110110011000",
    "1110111010101101",
    "1110111111000111",
    "1111000010101110",
    "1111000101000101",
    "1111000110010110",
    "1111000111011011",
    "1111001010100110",
    "1111010011000110",
    "1111100011001011",
    "1111111010110010",
    "1111101000111000",
    "1111001101000000",
    "1110110111001000",
    "1110101011101011",
    "1110101100011001",
    "1110110111100000",
    "1111001000111111",
    "1111011100011100",
    "1111101110011110",
    "1111111101011000",
    "1111110111000001",
    "1111101110010101",
    "1111100111110101",
    "1111100011010000",
    "1111100000111001",
    "1111100001000011",
    "1111100011101100",
    "1111101000000100",
    "1111101100101101",
    "1111110000000100",
    "1111110000111100",
    "1111101111000001",
    "1111101010101100",
    "1111100100111001",
    "1111011110101110",
    "1111011001011101",
    "1111010110000011",
    "1111010101010011",
    "1111010111100011",
    "1111011101000101",
    "1111100101111001",
    "1111110010000011",
    "1111111110100001",
    "1111101100010111",
    "1111011000011011",
    "1111000100010010",
    "1110110001100110",
    "1110100001110000",
    "1110010101101001",
    "1110001101100110",
    "1110001001110010",
    "1110001010100110",
    "1110010000100111",
    "1110011100010111",
    "1110101101101110",
    "1111000011101100",
    "1111011100001001",
    "1111110100010001",
    "1111110110110001",
    "1111100111011010",
    "1111011111000100",
    "1111011110000010",
    "1111100011110100",
    "1111101111000101",
    "1111111101111110",
    "1111110001101001",
    "1111100010001101",
    "1111010101110110",
    "1111001110001100",
    "1111001011110111",
    "1111001110011111",
    "1111010100110001",
    "1111011100111010",
    "1111100101001000",
    "1111101100000111",
    "1111110001011011",
    "1111110101010000",
    "1111111000010010",
    "1111111011010100",
    "1111111110111000",
    "1111111101000111",
    "1111111001011000",
    "1111110110111011",
    "1111110110101111",
    "1111111001011111",
    "1111111111011010",
    "1111110111100010",
    "1111101011100100",
    "1111011100101010",
    "1111001011000010",
    "1110110111110111",
    "1110100101010000",
    "1110010110010000",
    "1110001101110101",
    "1110001101111011",
    "1110010111000100",
    "1110101000000110",
    "1110111110111010",
    "1111011001010101",
    "1111110101100110",
    "1111101101111000",
    "1111010011000110",
    "1110111100010111",
    "1110101100001001",
    "1110100100010111",
    "1110100101110001",
    "1110101111110001",
    "1111000000011111",
    "1111010101101010",
    "1111101101010100",
    "1111111010000011",
    "1111100001111000",
    "1111001011100101",
    "1110111001000010",
    "1110101100001001",
    "1110100110000110",
    "1110100110111001",
    "1110101100110111",
    "1110110101000001",
    "1110111100001001",
    "1110111111101000",
    "1110111110011111",
    "1110111001100101",
    "1110110011000011",
    "1110101101011110",
    "1110101010110000",
    "1110101011100011",
    "1110101111010001",
    "1110110100101010",
    "1110111011000010",
    "1111000010111110",
    "1111001110000111",
    "1111011110001001",
    "1111110011011000",
    "1111110011101111",
    "1111011010101011",
    "1111000101100000",
    "1110110111100010",
    "1110110010000101",
    "1110110100000101",
    "1110111010110000",
    "1111000010111001",
    "1111001001110100",
    "1111001101111111",
    "1111001110111101",
    "1111001100111010",
    "1111001000011010",
    "1111000010000101",
    "1110111010101000",
    "1110110010111110",
    "1110101100001110",
    "1110100111011011",
    "1110100101100010",
    "1110100110101111",
    "1110101010100010",
    "1110110000000011",
    "1110110110101010",
    "1110111110011001",
    "1111001000000001",
    "1111010100101010",
    "1111100100111100",
    "1111111000010000",
    "1111110011001111",
    "1111100000011001",
    "1111010010000110",
    "1111001010011101",
    "1111001010000001",
    "1111001111110110",
    "1111011001111100",
    "1111100110000011",
    "1111110010001110",
    "1111111101001010",
    "1111111001111010",
    "1111110011110001",
    "1111110001000011",
    "1111110010011001",
    "1111111000000001",
    "1111111110011111",
    "1111110010100100",
    "1111100110000100",
    "1111011010110111",
    "1111010010001000",
    "1111001100000101",
    "1111001000001110",
    "1111000101101010",
    "1111000011110100",
    "1111000010011010",
    "1111000001101100",
    "1111000010000101",
    "1111000100001000",
    "1111001000000110",
    "1111001110001100",
    "1111010110011000",
    "1111100000100011",
    "1111101100010111",
    "1111111001010001",
    "1111111001011011",
    "1111101100101110",
    "1111100001100100",
    "1111011000101100",
    "1111010010100001",
    "1111001110110011",
    "1111001100111000",
    "1111001011101111",
    "1111001010010001",
    "1111000111111010",
    "1111000100101111",
    "1111000001011010",
    "1110111111000100",
    "1110111110110000",
    "1111000000111110",
    "1111000101010101",
    "1111001010100101",
    "1111001111000111",
    "1111010001010111",
    "1111010000011111",
    "1111001100100110",
    "1111000110111001",
    "1111000001010100",
    "1110111101111111",
    "1110111110111011",
    "1111000101110010",
    "1111010011110011",
    "1111101001000111",
    "1111111011110001",
    "1111011110001101",
    "1111000010100010",
    "1110101101000010",
    "1110100000101011",
    "1110011110010100",
    "1110100100011000",
    "1110101111100001",
    "1110111011110111",
    "1111000110010110",
    "1111001101010111",
    "1111010000110110",
    "1111010001110001",
    "1111010001011110",
    "1111010001000111",
    "1111010001010100",
    "1111010010000110",
    "1111010011001111",
    "1111010100011100",
    "1111010101101001",
    "1111010110111111",
    "1111011000101100",
    "1111011010101000",
    "1111011100110000",
    "1111011111000111",
    "1111100010001111",
    "1111100110110101",
    "1111101101101001",
    "1111110110110110",
    "1111111110000010",
    "1111110010001010",
    "1111100110110100",
    "1111011100111010",
    "1111010100011101",
    "1111001100101010",
    "1111000100001110",
    "1110111010010001",
    "1110101110101000",
    "1110100010001011",
    "1110010110011111",
    "1110001101001110",
    "1110000111011000",
    "1110000100111110",
    "1110000101000001",
    "1110000110001000",
    "1110000111000110",
    "1110000111011011",
    "1110001000011010",
    "1110001101000010",
    "1110011000010101",
    "1110101011011011",
    "1111000100100111",
    "1111011111011110",
    "1111110110011000",
    "1111111011110011",
    "1111111010000101",
    "1111111011111010",
    "1111101001001100",
    "1111010001101110",
    "1110111001100011",
    "1110100011111000",
    "1110010010110100",
    "1110000111101100",
    "1110000011000001",
    "1110000100110011",
    "1110001100101000",
    "1110011001101101",
    "1110101011001111",
    "1111000000110110",
    "1111011001111100",
    "1111110101010110",
    "1111101110111101",
    "1111010101110100",
    "1111000010001000",
    "1110110110010110",
    "1110110011101001",
    "1110111001010101",
    "1111000101001101",
    "1111010100101111",
    "1111100110000011",
    "1111111000010100",
    "1111110100011111",
    "1111100000110001",
    "1111001101100001",
    "1110111100101101",
    "1110110000100111",
    "1110101011000010",
    "1110101100101101",
    "1110110101000011",
    "1111000010011100",
    "1111010011000001",
    "1111100101001110",
    "1111110111110100",
    "1111110110011001",
    "1111100110110010",
    "1111011010111010",
    "1111010100001110",
    "1111010100000000",
    "1111011010110111",
    "1111101000100011",
    "1111111011110011",
    "1111101101100101",
    "1111010110101010",
    "1111000010010100",
    "1110110010111001",
    "1110101010001011",
    "1110101000110100",
    "1110101110011110",
    "1110111010000001",
    "1111001001110111",
    "1111011100100101",
    "1111110000111000",
    "1111111010011000",
    "1111100110011111",
    "1111010100101110",
    "1111000110001110",
    "1110111011111100",
    "1110110110011011",
    "1110110101110001",
    "1110111001100101",
    "1111000001001111",
    "1111001100001110",
    "1111011010010110",
    "1111101011100110",
    "1111111111011110",
    "1111101011100100",
    "1111010111111010",
    "1111001000001110",
    "1110111110101101",
    "1110111100100101",
    "1111000001110110",
    "1111001101100001",
    "1111011110011111",
    "1111110011111100",
    "1111110010110100",
    "1111010111000110",
    "1110111011010110",
    "1110100010111110",
    "1110010001100010",
    "1110001001110010",
    "1110001100111000",
    "1110011010011000",
    "1110110000011001",
    "1111001100001001",
    "1111101010000101",
    "1111111001100011",
    "1111100010001101",
    "1111010010100001",
    "1111001011110101",
    "1111001110010010",
    "1111011000111001",
    "1111101010000000",
    "1111111111110110",
    "1111100110010000",
    "1111001011000110",
    "1110110000111011",
    "1110011010101011",
    "1110001011000111",
    "1110000100000001",
    "1110000101110110",
    "1110001111101001",
    "1110011111011100",
    "1110110010110100",
    "1111000111101100",
    "1111011100100000",
    "1111110000010101",
    "1111111101010111",
    "1111101101010001",
    "1111100000000010",
    "1111010110010010",
    "1111010000010010",
    "1111001101110111",
    "1111001110011110",
    "1111010001011010",
    "1111010101111110",
    "1111011011101010",
    "1111100010000110",
    "1111101001010101",
    "1111110001110011",
    "1111111100011110",
    "1111110101100111",
    "1111100100001011",
    "1111010000010010",
    "1110111100011100",
    "1110101100000100",
    "1110100010000101",
    "1110011111110110",
    "1110100100101100",
    "1110101110010110",
    "1110111001110000",
    "1111000100100100",
    "1111001101111000",
    "1111010110100111",
    "1111100000011001",
    "1111101100101000",
    "1111111011011110",
    "1111110100100001",
    "1111100110001001",
    "1111011100010110",
    "1111011001010000",
    "1111011101010010",
    "1111100111011011",
    "1111110101100100",
    "1111111010011010",
    "1111101010011010",
    "1111011011101000",
    "1111001111000111",
    "1111000110000000",
    "1111000001100010",
    "1111000010110100",
    "1111001010011000",
    "1111010111100010",
    "1111101000100100",
    "1111111010101101",
    "1111110100111011",
    "1111101000101010",
    "1111100001011111",
    "1111011111001000",
    "1111100000011111",
    "1111100100001011",
    "1111101001000101",
    "1111101110100110",
    "1111110100100100",
    "1111111011001000",
    "1111111101100000",
    "1111110101010100",
    "1111101100011101",
    "1111100011011010",
    "1111011011000001",
    "1111010100011000",
    "1111010000110110",
    "1111010001100010",
    "1111010111000001",
    "1111100001000101",
    "1111101110100111",
    "1111111101111010",
    "1111110011000001",
    "1111100110010000",
    "1111011101011110",
    "1111011010000001",
    "1111011100111101",
    "1111100110110011",
    "1111110111001010",
    "1111110011011111",
    "1111011011111000",
    "1111000101000101",
    "1110110010000000",
    "1110100100100101",
    "1110011101011110",
    "1110011100000101",
    "1110011111000101",
    "1110100100110111",
    "1110101100010011",
    "1110110100101110",
    "1110111110001010",
    "1111001001000001",
    "1111010101101100",
    "1111100100001101",
    "1111110100000010",
    "1111111011111111",
    "1111101101101100",
    "1111100010111101",
    "1111011101101000",
    "1111011111010001",
    "1111101000111100",
    "1111111010100010",
    "1111101101101010",
    "1111010010111011",
    "1110111001010001",
    "1110100100101010",
    "1110010111111001",
    "1110010100000110",
    "1110011000011010",
    "1110100010100001",
    "1110101111111101",
    "1110111111100100",
    "1111010001100111",
    "1111100110111000",
    "1111111111000111",
    "1111100111101010",
    "1111010001010101",
    "1111000010011010",
    "1110111110110001",
    "1111001000100101",
    "1111011111011010",
    "1111111111110100",
    "1111011010010100",
    "1110110101110110",
    "1110010111011010",
    "1110000010100100",
    "1101111000110101",
    "1101111001100011",
    "1110000010001101",
    "1110001111011100",
    "1110011110001010",
    "1110101100010001",
    "1110111001001011",
    "1111000101100000",
    "1111010010111000",
    "1111100011001000",
    "1111110111011011",
    "1111110000011011",
    "1111010110001011",
    "1110111100100001",
    "1110100110010101",
    "1110010101101100",
    "1110001011011001",
    "1110000110111111",
    "1110000111010101",
    "1110001011000001",
    "1110010000100100",
    "1110010110110010",
    "1110011100101011",
    "1110100001011111",
    "1110100100100100",
    "1110100101100101",
    "1110100101010111",
    "1110100110011000",
    "1110101011110111",
    "1110111000000110",
    "1111001011001110",
    "1111100010101011",
    "1111111001110100",
    "1111110100010111",
    "1111101011100101",
    "1111101100010111",
    "1111110100010101",
    "1111111111100110",
    "1111110101011010",
    "1111101100110101",
    "1111100110101010",
    "1111100001101011",
    "1111011100010001",
    "1111010101110001",
    "1111001110111010",
    "1111001001100010",
    "1111000111110001",
    "1111001010111100",
    "1111010010111000",
    "1111011101101011",
    "1111101000100111",
    "1111110001001010",
    "1111110101100110",
    "1111110101011101",
    "1111110001011000",
    "1111101011000011",
    "1111100100101001",
    "1111100000010010",
    "1111011111011001",
    "1111100010100001",
    "1111101001001101",
    "1111110010010101",
    "1111111100010110",
    "1111111010001010",
    "1111110010010010",
    "1111101100010110",
    "1111101000000010",
    "1111100100101010",
    "1111100001010000",
    "1111011101001110",
    "1111011000011011",
    "1111010011101001",
    "1111010000000011",
    "1111001111001010",
    "1111010010001111",
    "1111011010000111",
    "1111100111001111",
    "1111111001010100",
    "1111110000101101",
    "1111011000110000",
    "1111000001010101",
    "1110101101001100",
    "1110011110101101",
    "1110010111010011",
    "1110010111010101",
    "1110011101111101",
    "1110101001010110",
    "1110110111010000",
    "1111000101010011",
    "1111010001011010",
    "1111011010000010",
    "1111011110010100",
    "1111011110000101",
    "1111011001111001",
    "1111010010111011",
    "1111001010100010",
    "1111000010000010",
    "1110111010011000",
    "1110110100001000",
    "1110101111011100",
    "1110101100010100",
    "1110101010110111",
    "1110101011010110",
    "1110101110001100",
    "1110110011110011",
    "1110111100100001",
    "1111001000110100",
    "1111011001000110",
    "1111101101101000",
    "1111111001111101",
    "1111011111100011",
    "1111000110000110",
    "1110110001010000",
    "1110100100001000",
    "1110100000011110",
    "1110100110000000",
    "1110110010110011",
    "1111000100000001",
    "1111010111010000",
    "1111101011010111",
    "1111111111010011",
    "1111101000000011",
    "1111001110101000",
    "1110110100011000",
    "1110011100010110",
    "1110001010011101",
    "1110000010001011",
    "1110000101010011",
    "1110010011000110",
    "1110101000101010",
    "1111000001110110",
    "1111011010011011",
    "1111101110111110",
    "1111111101010111",
    "1111111011001100",
    "1111111010011101",
    "1111111111001100",
    "1111111000010010",
    "1111101110001011",
    "1111100100101001",
    "1111011101110000",
    "1111011011100000",
    "1111011111001000",
    "1111101000111010",
    "1111110111100011",
    "1111110111011100",
    "1111100111011101",
    "1111011011100101",
    "1111010110000100",
    "1111011000001000",
    "1111100001101100",
    "1111110001100011",
    "1111111010100011",
    "1111100101100101",
    "1111010010011101",
    "1111000011100111",
    "1110111010011110",
    "1110110111001110",
    "1110111001000010",
    "1110111110110001",
    "1111000111110100",
    "1111010100011010",
    "1111100101000110",
    "1111111001111101",
    "1111101110001111",
    "1111010110000110",
    "1111000000101011",
    "1110110000101001",
    "1110100111001110",
    "1110100011111011",
    "1110100100110001",
    "1110100111011111",
    "1110101010100110",
    "1110101110010110",
    "1110110100000110",
    "1110111101011110",
    "1111001010110111",
    "1111011010110010",
    "1111101010001110",
    "1111110101010001",
    "1111111000100110",
    "1111110010101100",
    "1111100100011010",
    "1111010000110011",
    "1110111100000101",
    "1110101010011011",
    "1110011111000100",
    "1110011011110010",
    "1110100001000111",
    "1110101110010111",
    "1111000010010010",
    "1111011010111101",
    "1111110110001000",
    "1111101110110111",
    "1111010110111001",
    "1111000100010111",
    "1110111000110010",
    "1110110100100100",
    "1110110110111011",
    "1110111110010111",
    "1111001001011000",
    "1111010110110010",
    "1111100110000000",
    "1111110110100110",
    "1111110111110101",
    "1111100110000001",
    "1111010100111110",
    "1111000101110010",
    "1110111001100010",
    "1110110000110101",
    "1110101100000100",
    "1110101011100101",
    "1110101111100011",
    "1110111000001011",
    "1111000101001000",
    "1111010101010111",
    "1111100110110010",
    "1111110110101001",
    "1111111110000001",
    "1111111001101011",
    "1111111101010101",
    "1111110111101110",
    "1111100111111000",
    "1111010110010000",
    "1111000110001000",
    "1110111010000110",
    "1110110011101111",
    "1110110011100010",
    "1110111001000110",
    "1111000011011111",
    "1111010001110000",
    "1111100011000001",
    "1111110110101000",
    "1111110011111110",
    "1111011101100011",
    "1111000111010101",
    "1110110011001010",
    "1110100011001101",
    "1110011001100011",
    "1110010111011000",
    "1110011100101101",
    "1110101000001011",
    "1110110111011000",
    "1111000111011101",
    "1111010110000001",
    "1111100001101100",
    "1111101011001001",
    "1111110100111101",
    "1111111110000111",
    "1111101100110111",
    "1111011000101100",
    "1111000101011111",
    "1110111000011000",
    "1110110110000110",
    "1111000001000101",
    "1111011000010000",
    "1111110111011110",
    "1111100111000110",
    "1111001001011000",
    "1110110011100111",
    "1110101000000011",
    "1110100110101010",
    "1110101101110000",
    "1110111010110000",
    "1111001010111111",
    "1111011100000100",
    "1111101011111001",
    "1111111000110000",
    "1111111110110111",
    "1111111100000011",
    "1111111110111011",
    "1111111001100000",
    "1111101111001110",
    "1111100100101001",
    "1111011100000101",
    "1111010111100010",
    "1111010111111110",
    "1111011101010010",
    "1111100110010011",
    "1111110000110110",
    "1111111010011001",
    "1111111111001100",
    "1111111101011010",
    "1111111111100101",
    "1111111000111110",
    "1111110000110010",
    "1111101001100001",
    "1111100101010101",
    "1111100101100111",
    "1111101010111000",
    "1111110100110011",
    "1111111101011000",
    "1111101100110010",
    "1111011010111000",
    "1111001001100000",
    "1110111010110101",
    "1110110000110000",
    "1110101100100011",
    "1110101110010100",
    "1110110101000001",
    "1110111110110001",
    "1111001001111001",
    "1111010101110001",
    "1111100010111001",
    "1111110010010110",
    "1111111011011100",
    "1111100111011000",
    "1111010011100001",
    "1111000010101100",
    "1110110111101000",
    "1110110011110011",
    "1110110111000001",
    "1111000000000000",
    "1111001101001010",
    "1111011101111000",
    "1111110010010101",
    "1111110101000111",
    "1111011001000110",
    "1110111011111100",
    "1110100001011111",
    "1110001110010010",
    "1110000110010011",
    "1110001011011110",
    "1110011100111111",
    "1110110111011010",
    "1111010101100010",
    "1111110001111001",
    "1111110111111100",
    "1111101010100011",
    "1111100110011100",
    "1111101010011110",
    "1111110100101010",
    "1111111100110101",
    "1111101011101010",
    "1111011001000100",
    "1111000110100000",
    "1110110101101010",
    "1110101000001110",
    "1110011111010001",
    "1110011011001010",
    "1110011011100110",
    "1110011111110101",
    "1110100111010101",
    "1110110010010101",
    "1111000001101011",
    "1111010110001001",
    "1111101111101000",
    "1111110011101000",
    "1111010111000011",
    "1110111110101011",
    "1110101110010010",
    "1110101000000011",
    "1110101100001111",
    "1110111001100011",
    "1111001101111111",
    "1111100111100101",
    "1111111011011001",
    "1111011100111111",
    "1110111111101000",
    "1110100110001101",
    "1110010011100111",
    "1110001001101101",
    "1110001000110100",
    "1110001111101001",
    "1110011100000010",
    "1110101011100101",
    "1110111100101000",
    "1111001110101101",
    "1111100010001101",
    "1111110111101101",
    "1111110001000010",
    "1111011001111001",
    "1111000101100111",
    "1110110111001011",
    "1110110000010101",
    "1110110001000010",
    "1110110111011010",
    "1111000000101001",
    "1111001010000111",
    "1111010010100110",
    "1111011010001110",
    "1111100010000000",
    "1111101010101010",
    "1111110011101100",
    "1111111011001100",
    "1111111110100111",
    "1111111011101001",
    "1111110001100111",
    "1111100001111001",
    "1111001111101100",
    "1110111111000010",
    "1110110011100010",
    "1110101111011111",
    "1110110011111100",
    "1111000001001010",
    "1111010110111011",
    "1111110100000100",
    "1111101010000011",
    "1111000111101101",
    "1110101001101010",
    "1110010100000101",
    "1110001001011011",
    "1110001001100010",
    "1110010001110100",
    "1110011110010001",
    "1110101010110101",
    "1110110101000000",
    "1110111011111111",
    "1111000000110110",
    "1111000101110001",
    "1111001101010100",
    "1111011001011000",
    "1111101010100001",
    "1111111111100111",
    "1111101001011010",
    "1111010011011010",
    "1111000000111101",
    "1110110011111001",
    "1110101100111000",
    "1110101011011011",
    "1110101110001001",
    "1110110011011100",
    "1110111010000111",
    "1111000010001111",
    "1111001100111000",
    "1111011011100011",
    "1111101110111100",
    "1111111001111010",
    "1111100001111000",
    "1111001100100000",
    "1110111100111111",
    "1110110100111110",
    "1110110100000101",
    "1110111000010000",
    "1110111110111101",
    "1111000110011011",
    "1111001110011110",
    "1111011000010101",
    "1111100101101001",
    "1111110111011110",
    "1111110010111011",
    "1111011100010001",
    "1111001000010001",
    "1110111010110000",
    "1110110110001110",
    "1110111011101101",
    "1111001010110100",
    "1111100001110110",
    "1111111101111010",
    "1111100100110100",
    "1111001010100101",
    "1110110111001000",
    "1110101100110111",
    "1110101100010111",
    "1110110100001011",
    "1111000001010100",
    "1111010000100100",
    "1111011111100110",
    "1111101101010101",
    "1111111001110000",
    "1111111011000000",
    "1111110001010110",
    "1111101010011111",
    "1111101000010000",
    "1111101100010011",
    "1111110111001011",
    "1111111000001011",
    "1111100100011000",
    "1111010000100100",
    "1110111111100001",
    "1110110010101111",
    "1110101010100101",
    "1110100110100000",
    "1110100101111001",
    "1110101000010110",
    "1110101101110101",
    "1110110110011011",
    "1111000010010010",
    "1111010001100010",
    "1111100100010010",
    "1111111010011001",
    "1111101100111011",
    "1111010011011100",
    "1110111011101101",
    "1110101000110100",
    "1110011101100001",
    "1110011011101010",
    "1110100011000110",
    "1110110001110100",
    "1111000100010101",
    "1111010110100101",
    "1111100101001000",
    "1111101101101110",
    "1111101111110010",
    "1111101011111100",
    "1111100011100100",
    "1111011000001110",
    "1111001011001100",
    "1110111101101001",
    "1110110000011110",
    "1110100100010101",
    "1110011001110000",
    "1110010001000101",
    "1110001010011011",
    "1110000101111100",
    "1110000011101110",
    "1110000011111100",
    "1110000110111100",
    "1110001101100100",
    "1110011001010001",
    "1110101011001110",
    "1111000011010111",
    "1111011111101011",
    "1111111100001100",
    "1111101011110111",
    "1111011100110010",
    "1111011000111001",
    "1111011111111000",
    "1111101111100000",
    "1111111011000001",
    "1111100001110100",
    "1111000101111110",
    "1110101000011101",
    "1110001011000111",
    "1101110000111011",
    "1101011101011100",
    "1101010011110110",
    "1101010101100100",
    "1101100001011100",
    "1101110100000101",
    "1110001001001001",
    "1110011101111011",
    "1110110010011101",
    "1111001000100011",
    "1111100010000000",
    "1111111110101000",
    "1111100100011000",
    "1111001011110000",
    "1110111100001111",
    "1110111000100101",
    "1111000000001000",
    "1111001111100011",
    "1111100010010010",
    "1111110100011010",
    "1111111011110011",
    "1111101110010100",
    "1111100001110110",
    "1111010101000101",
    "1111000111101010",
    "1110111010100011",
    "1110101111010110",
    "1110100111100011",
    "1110100011111100",
    "1110100100000101",
    "1110100110101100",
    "1110101010100101",
    "1110101111000000",
    "1110110011111001",
    "1110111001100000",
    "1111000000010111",
    "1111001001001011",
    "1111010100100111",
    "1111100010111011",
    "1111110011100110",
    "1111111010110011",
    "1111101010100101",
    "1111011110000000",
    "1111010110101101",
    "1111010101000110",
    "1111011000001110",
    "1111011110001010",
    "1111100100110100",
    "1111101010100010",
    "1111101110101010",
    "1111110001100010",
    "1111110100000010",
    "1111110110111111",
    "1111111010100100",
    "1111111110000011",
    "1111111111110110",
    "1111111111011000",
    "1111111011010001",
    "1111110100001100",
    "1111101011011100",
    "1111100010101001",
    "1111011011011001",
    "1111010110111110",
    "1111010110010010",
    "1111011001110000",
    "1111100001010111",
    "1111101100100101",
    "1111111010100011",
    "1111110101111000",
    "1111100110001110",
    "1111011000000011",
    "1111001100110000",
    "1111000101100100",
    "1111000011000101",
    "1111000101011011",
    "1111001100000101",
    "1111010110000100",
    "1111100010000011",
    "1111101110110011",
    "1111111011001001",
    "1111111001101001",
    "1111110000001000",
    "1111101000011011",
    "1111100010100010",
    "1111011110011100",
    "1111011100001110",
    "1111011011111100",
    "1111011101101110",
    "1111100001011110",
    "1111100110100100",
    "1111101100000100",
    "1111110000101111",
    "1111110011001110",
    "1111110010010001",
    "1111101101001000",
    "1111100011111000",
    "1111010111101010",
    "1111001010010110",
    "1110111110001001",
    "1110110100111011",
    "1110101111111010",
    "1110101111100001",
    "1110110011011010",
    "1110111010110101",
    "1111000100111100",
    "1111010001000101",
    "1111011110100011",
    "1111101100100011",
    "1111111010000110",
    "1111111001111101",
    "1111110000110110",
    "1111101011010100",
    "1111101001101000",
    "1111101011010001",
    "1111101111010001",
    "1111110100011111",
    "1111111010000110",
    "1111111111110000",
    "1111111010000111",
    "1111110010110010",
    "1111101001000110",
    "1111011100000101",
    "1111001011001110",
    "1110110111000100",
    "1110100001100111",
    "1110001101110101",
    "1101111110111011",
    "1101110111010101",
    "1101110111110100",
    "1101111111011110",
    "1110001100000100",
    "1110011011000100",
    "1110101010100010",
    "1110111001110010",
    "1111001000111001",
    "1111010111111110",
    "1111100110010011",
    "1111110010010100",
    "1111111001110000",
    "1111111010100100",
    "1111110011110000",
    "1111100110000001",
    "1111010011101100",
    "1111000000000000",
    "1110101110001010",
    "1110100000100011",
    "1110011000010000",
    "1110010101000011",
    "1110010101110111",
    "1110011001001011",
    "1110011101011001",
    "1110100001010100",
    "1110100100010010",
    "1110100110011010",
    "1110101000011010",
    "1110101011011101",
    "1110110000111000",
    "1110111001111001",
    "1111000111001110",
    "1111011000110101",
    "1111101101100101",
    "1111111100101100",
    "1111101000101111",
    "1111011000111111",
    "1111001111000010",
    "1111001011001100",
    "1111001100100001",
    "1111010001000011",
    "1111010110100000",
    "1111011010111010",
    "1111011101001010",
    "1111011101010010",
    "1111011100111111",
    "1111011110110110",
    "1111100101010011",
    "1111110001010010",
    "1111111110011011",
    "1111101101000010",
    "1111011110100001",
    "1111010110011101",
    "1111010110101000",
    "1111011110100100",
    "1111101100000110",
    "1111111100100000",
    "1111110010100100",
    "1111100010111011",
    "1111010101101110",
    "1111001100000100",
    "1111000110111110",
    "1111000111100101",
    "1111001110110001",
    "1111011100110010",
    "1111110000111111",
    "1111110110001010",
    "1111011011011011",
    "1111000010001010",
    "1110101101101011",
    "1110100000011111",
    "1110011011111000",
    "1110011111101011",
    "1110101010011000",
    "1110111001100011",
    "1111001010100010",
    "1111011010111000",
    "1111101001000000",
    "1111110011111011",
    "1111111011010101",
    "1111111111001111",
    "1111111111111000",
    "1111111101100001",
    "1111111000100110",
    "1111110001100111",
    "1111101001001100",
    "1111100000000011",
    "1111010110110100",
    "1111001101111011",
    "1111000101101010",
    "1110111110001111",
    "1110110111111001",
    "1110110010111110",
    "1110101111110001",
    "1110101110101110",
    "1110110000011001",
    "1110110101100000",
    "1110111110110101",
    "1111001100100110",
    "1111011110001001",
    "1111110001101000",
    "1111111011100101",
    "1111101100010111",
    "1111100010110110",
    "1111011111110000",
    "1111100010001011",
    "1111101000000100",
    "1111101110101110",
    "1111110011111000",
    "1111110110000101",
    "1111110101000111",
    "1111110001100110",
    "1111101100101100",
    "1111100111011000",
    "1111100010000010",
    "1111011100000100",
    "1111010100011010",
    "1111001001110101",
    "1110111011110000",
    "1110101010100010",
    "1110010111110001",
    "1110000110000000",
    "1101111000000100",
    "1101110000001111",
    "1101101111011100",
    "1101110101000011",
    "1101111111001000",
    "1110001011001111",
    "1110010111000100",
    "1110100001000011",
    "1110101001110101",
    "1110110100111001",
    "1111000101111011",
    "1111011110010111",
    "1111111100000011",
    "1111100110011101",
    "1111001111110000",
    "1111000100111011",
    "1111001000001000",
    "1111010110110110",
    "1111101011100011",
    "1111111111101011",
    "1111101111010110",
    "1111100101000001",
    "1111100000010001",
    "1111011111110110",
    "1111100010100111",
    "1111100111110110",
    "1111101111011101",
    "1111111001001010",
    "1111111011111100",
    "1111110001011101",
    "1111101001011000",
    "1111100101011000",
    "1111100101111110",
    "1111101010001010",
    "1111110000001000",
    "1111110110001000",
    "1111111011001101",
    "1111111111000111",
    "1111111101110111",
    "1111111011001000",
    "1111110111101110",
    "1111110010100011",
    "1111101010011000",
    "1111011110001001",
    "1111001101101000",
    "1110111001101011",
    "1110100100101001",
    "1110010001100110",
    "1110000011101111",
    "1101111101010100",
    "1101111110111010",
    "1110000111001011",
    "1110010011010011",
    "1110011111111000",
    "1110101001110111",
    "1110101111101000",
    "1110110001010101",
    "1110110001011110",
    "1110110011110001",
    "1110111011011011",
    "1111001001100010",
    "1111011100100110",
    "1111110001000011",
    "1111111101011010",
    "1111110010100111",
    "1111110000011101",
    "1111110110010100",
    "1111111110000011",
    "1111101111001110",
    "1111011111001010",
    "1111001111001111",
    "1111000000110101",
    "1110110101101001",
    "1110101111110000",
    "1110110001100010",
    "1110111100111101",
    "1111010010011100",
    "1111101111111010",
    "1111101110110100",
    "1111001111001111",
    "1110110110000100",
    "1110100110010000",
    "1110100000001101",
    "1110100010010010",
    "1110101001111101",
    "1110110101001011",
    "1111000010110011",
    "1111010010100001",
    "1111100100001110",
    "1111110111001011",
    "1111110110010010",
    "1111100110011011",
    "1111011011011001",
    "1111010110100000",
    "1111011000000011",
    "1111011111001100",
    "1111101010011111",
    "1111111000000001",
    "1111111001111011",
    "1111101100110110",
    "1111100001110000",
    "1111011001011000",
    "1111010100011000",
    "1111010011011000",
    "1111010110110100",
    "1111011111001111",
    "1111101101011010",
    "1111111110001011",
    "1111100100001011",
    "1111000110101100",
    "1110101001001011",
    "1110001111101001",
    "1101111101110101",
    "1101110101110001",
    "1101110111011111",
    "1110000000110110",
    "1110001110101011",
    "1110011101110111",
    "1110101100111100",
    "1110111100101011",
    "1111001111011001",
    "1111100111000101",
    "1111111100000000",
    "1111011100100001",
    "1110111111000101",
    "1110101000101111",
    "1110011101000101",
    "1110011100101101",
    "1110100101001011",
    "1110110010010000",
    "1110111111111000",
    "1111001100001111",
    "1111011000001100",
    "1111100110001101",
    "1111111000010111",
    "1111110001001011",
    "1111011001010000",
    "1111000100101100",
    "1110111000101111",
    "1110111001001110",
    "1111000111001000",
    "1111100000100100",
    "1111111110011011",
    "1111011011000111",
    "1110111010101101",
    "1110100001011111",
    "1110010010011010",
    "1110001110100100",
    "1110010101011101",
    "1110100101010000",
    "1110111011011000",
    "1111010101010011",
    "1111110000111000",
    "1111110011111110",
    "1111011011110010",
    "1111001000111110",
    "1110111101110111",
    "1110111100010001",
    "1111000101001000",
    "1111011000001000",
    "1111110011001100",
    "1111101101011000",
    "1111001110010010",
    "1110110100001000",
    "1110100010000010",
    "1110011001000001",
    "1110011000000011",
    "1110011100101010",
    "1110100100010010",
    "1110101101001100",
    "1110110110111011",
    "1111000010000110",
    "1111001111110101",
    "1111100000111011",
    "1111110101100001",
    "1111110011010100",
    "1111011011101000",
    "1111000101110001",
    "1110110011111110",
    "1110100111100000",
    "1110100000101011",
    "1110011110111010",
    "1110100001100010",
    "1110100111110111",
    "1110110001100001",
    "1110111110011111",
    "1111001110111111",
    "1111100011000001",
    "1111111010000011",
    "1111101101100110",
    "1111010110101000",
    "1111000011111110",
    "1110110111110101",
    "1110110010111101",
    "1110110100010011",
    "1110111001100011",
    "1111000000000000",
    "1111000101101001",
    "1111001001110101",
    "1111001101100011",
    "1111010010101011",
    "1111011011010011",
    "1111101000100001",
    "1111111010000000",
    "1111110010000111",
    "1111011111000100",
    "1111010000000000",
    "1111000111011000",
    "1111000110001001",
    "1111001011101010",
    "1111010110010101",
    "1111100100010000",
    "1111110011011110",
    "1111111101111001",
    "1111110001111100",
    "1111101010101111",
    "1111101010000111",
    "1111110001001000",
    "1111111111100001",
    "1111101100101000",
    "1111010110101100",
    "1111000010101011",
    "1110110100001110",
    "1110101101100001",
    "1110101110110000",
    "1110110110001101",
    "1111000001000101",
    "1111001100100001",
    "1111010110101000",
    "1111011111011001",
    "1111101000101011",
    "1111110101001011",
    "1111111001001000",
    "1111100010010010",
    "1111001000100010",
    "1110101111111111",
    "1110011101000101",
    "1110010011011010",
    "1110010100010010",
    "1110011110101110",
    "1110110000011001",
    "1111000110100111",
    "1111011111001111",
    "1111111000101001",
    "1111101110011000",
    "1111010111010011",
    "1111000011101110",
    "1110110101011101",
    "1110101110000101",
    "1110101110001010",
    "1110110101001101",
    "1111000001010100",
    "1111001111111010",
    "1111011110001101",
    "1111101010000110",
    "1111110010010011",
    "1111110110101010",
    "1111110111110011",
    "1111110110110011",
    "1111110100111011",
    "1111110011001001",
    "1111110001111011",
    "1111110001001100",
    "1111110000011011",
    "1111101110111100",
    "1111101100010010",
    "1111101000011001",
    "1111100011111001",
    "1111100000000010",
    "1111011110010111",
    "1111100000011111",
    "1111100111101011",
    "1111110100100111",
    "1111111000101001",
    "1111100001001000",
    "1111000110111001",
    "1110101100111111",
    "1110010110111111",
    "1110001000010011",
    "1110000011011101",
    "1110001001111001",
    "1110011011100101",
    "1110110110111001",
    "1111011000100010",
    "1111111100000011",
    "1111100011011010",
    "1111001010000111",
    "1110111010110000",
    "1110110110001000",
    "1110111011000100",
    "1111000111010101",
    "1111011000111110",
    "1111101111000111",
    "1111110110010100",
    "1111010111110100",
    "1110110111001001",
    "1110010111100010",
    "1101111100110011",
    "1101101010010110",
    "1101100001110110",
    "1101100010110001",
    "1101101010110000",
    "1101110110100111",
    "1110000011100010",
    "1110010000000000",
    "1110011011100110",
    "1110100110100100",
    "1110110001001000",
    "1110111011000111",
    "1111000100001010",
    "1111001011110111",
    "1111010010010010",
    "1111011000001011",
    "1111011110101101",
    "1111100110110111",
    "1111110000111101",
    "1111111100011100",
    "1111110111110011",
    "1111101100111110",
    "1111100011110100",
    "1111011100100000",
    "1111010110110111",
    "1111010010110110",
    "1111010000100100",
    "1111010000100100",
    "1111010011101110",
    "1111011010110100",
    "1111100110000110",
    "1111110100111100",
    "1111111010001111",
    "1111101001101110",
    "1111011011100110",
    "1111010001011010",
    "1111001011110111",
    "1111001010110101",
    "1111001101110011",
    "1111010100000101",
    "1111011101000100",
    "1111100111110011",
    "1111110010110101",
    "1111111100000011",
    "1111111110110001",
    "1111111111101111",
    "1111110111111011",
    "1111101000010001",
    "1111010010110100",
    "1110111010100110",
    "1110100011011000",
    "1110010000101100",
    "1110000101000101",
    "1110000001100001",
    "1110000101011111",
    "1110001111011111",
    "1110011101111111",
    "1110101111111111",
    "1111000101001000",
    "1111011101010100",
    "1111110111111111",
    "1111101100011000",
    "1111010010011010",
    "1110111100111101",
    "1110101110011100",
    "1110101000000011",
    "1110101001011011",
    "1110110001000000",
    "1110111100100110",
    "1111001010010001",
    "1111011000101100",
    "1111100111001101",
    "1111110101100010",
    "1111111100110011",
    "1111110000101001",
    "1111100110111111",
    "1111100000110011",
    "1111011110110000",
    "1111100000111101",
    "1111100110111000",
    "1111101111011110",
    "1111111001010101",
    "1111111100111101",
    "1111110100101000",
    "1111101110100011",
    "1111101011001001",
    "1111101010010101",
    "1111101011101000",
    "1111101110001110",
    "1111110001001000",
    "1111110011010001",
    "1111110011110111",
    "1111110010011011",
    "1111101111000010",
    "1111101010000010",
    "1111100100000001",
    "1111011101100110",
    "1111010111000011",
    "1111010000011110",
    "1111001001101011",
    "1111000010100100",
    "1110111011001100",
    "1110110011111001",
    "1110101101010010",
    "1110101000010000",
    "1110100101100111",
    "1110100110001011",
    "1110101010101010",
    "1110110011111000",
    "1111000010101111",
    "1111010111111110",
    "1111110011010010",
    "1111101101010011",
    "1111001101101011",
    "1110110010011100",
    "1110011111110001",
    "1110011000001000",
    "1110011011010100",
    "1110100110110110",
    "1110110110101100",
    "1111000111000100",
    "1111010101101010",
    "1111100010010000",
    "1111101101111001",
    "1111111001110011",
    "1111111001111110",
    "1111101111000101",
    "1111101000000111",
    "1111100111100100",
    "1111101110100001",
    "1111111011110100",
    "1111110011100101",
    "1111100011110001",
    "1111011000000110",
    "1111010010100001",
    "1111010011000110",
    "1111011000101100",
    "1111100001010101",
    "1111101011001100",
    "1111110100101010",
    "1111111100100011",
    "1111111101110001",
    "1111111010110100",
    "1111111010100111",
    "1111111100111110",
    "1111111110101101",
    "1111111001100000",
    "1111110100101011",
    "1111110001100010",
    "1111110001010001",
    "1111110100111011",
    "1111111101001001",
    "1111110110001110",
    "1111100110011100",
    "1111010101011111",
    "1111000101111001",
    "1110111010000001",
    "1110110011110100",
    "1110110100011111",
    "1110111100010110",
    "1111001010100011",
    "1111011101000000",
    "1111110000011101",
    "1111111110101111",
    "1111110011111111",
    "1111110001001101",
    "1111110110010110",
    "1111111110100011",
    "1111110000110101",
    "1111100011111011",
    "1111011010011000",
    "1111010101010011",
    "1111010100011111",
    "1111010110000100",
    "1111010110101010",
    "1111010010110001",
    "1111001000100000",
    "1110111000100011",
    "1110100110010110",
    "1110010110111100",
    "1110001111011001",
    "1110010011100010",
    "1110100100010111",
    "1110111111110000",
    "1111100001001111",
    "1111111101000101",
    "1111100000110001",
    "1111001101110111",
    "1111000110010011",
    "1111001001111100",
    "1111010111001001",
    "1111101011100110",
    "1111111011001000",
    "1111011111100011",
    "1111000100000001",
    "1110101011000100",
    "1110010110111011",
    "1110001000111111",
    "1110000001100100",
    "1101111111101001",
    "1110000001100001",
    "1110000101001001",
    "1110001000110111",
    "1110001011011101",
    "1110001100100011",
    "1110001100011110",
    "1110001100001001",
    "1110001100100000",
    "1110001110001010",
    "1110010001001000",
    "1110010100111001",
    "1110011000100111",
    "1110011011001111",
    "1110011011111101",
    "1110011010001110",
    "1110010101111100",
    "1110001111110000",
    "1110001000111111",
    "1110000100011010",
    "1110000101111001",
    "1110010001000011",
    "1110100111011111",
    "1111000111111001",
    "1111101110000100",
    "1111101011110110",
    "1111001011111100",
    "1110110110011101",
    "1110101100101101",
    "1110101100110111",
    "1110110011010111",
    "1110111100011100",
    "1111000101011010",
    "1111001101001010",
    "1111010011111100",
    "1111011011000111",
    "1111100100100000",
    "1111110001011111",
    "1111111101101101",
    "1111101010011111",
    "1111010111011111",
    "1111000111110010",
    "1110111101110011",
    "1110111010110000",
    "1110111110010100",
    "1111000111001101",
    "1111010011111100",
    "1111100011101100",
    "1111110110011011",
    "1111110011110100",
    "1111011100000111",
    "1111000100110110",
    "1110110001011100",
    "1110100101011000",
    "1110100010111011",
    "1110101010001111",
    "1110111001100000",
    "1111001101011110",
    "1111100010011101",
    "1111110101001111",
    "1111111100100101",
    "1111110100100100",
    "1111110011011111",
    "1111111001011100",
    "1111111010001101",
    "1111101001001011",
    "1111010101110111",
    "1111000011001111",
    "1110110011111011",
    "1110101001110101",
    "1110100101101100",
    "1110100110110100",
    "1110101011010110",
    "1110110000111000",
    "1110110101001000",
    "1110110110100101",
    "1110110100110111",
    "1110110000101100",
    "1110101011100110",
    "1110100111011011",
    "1110100101111100",
    "1110101000011010",
    "1110101111101100",
    "1110111100011110",
    "1111001110110110",
    "1111100101111100",
    "1111111111010101",
    "1111101000101001",
    "1111010101110111",
    "1111001011001010",
    "1111001001100000",
    "1111001111100100",
    "1111011010010100",
    "1111100110010000",
    "1111110001000001",
    "1111111010100101",
    "1111111010111110",
    "1111101101010001",
    "1111011011000110",
    "1111000101100100",
    "1110110000001101",
    "1110011111100001",
    "1110010111011111",
    "1110011010000001",
    "1110100110100101",
    "1110111011000111",
    "1111010101001000",
    "1111110010011111",
    "1111101110101111",
    "1111010000110110",
    "1110110110100101",
    "1110100010110001",
    "1110010111110001",
    "1110010110101000",
    "1110011110101001",
    "1110101101100110",
    "1111000000110101",
    "1111010101111001",
    "1111101011010010",
    "1111111111111011",
    "1111101100101010",
    "1111011100001111",
    "1111010000110001",
    "1111001100011110",
    "1111010000101110",
    "1111011100111111",
    "1111101110110000",
    "1111111101111011",
    "1111101101001100",
    "1111100001111101",
    "1111011101010010",
    "1111011110110110",
    "1111100101100101",
    "1111110000111101",
    "1111111110111100",
    "1111101010000111",
    "1111010001011010",
    "1110110111000011",
    "1110011110000100",
    "1110001001101111",
    "1101111100011011",
    "1101110110110111",
    "1101111000000001",
    "1101111101101000",
    "1110000101011111",
    "1110001110101110",
    "1110011010010001",
    "1110101010010110",
    "1111000000110000",
    "1111011101011001",
    "1111111101101010",
    "1111100010111101",
    "1111001001101011",
    "1110111010100010",
    "1110110111001011",
    "1110111110010010",
    "1111001100010111",
    "1111011101001010",
    "1111101101001011",
    "1111111010010010",
    "1111111100001000",
    "1111110101100101",
    "1111110000111100",
    "1111101101010001",
    "1111101010010001",
    "1111101000011000",
    "1111101000011010",
    "1111101011010110",
    "1111110001111000",
    "1111111100000111",
    "1111110110011110",
    "1111100111010101",
    "1111011000011110",
    "1111001100011011",
    "1111000101010000",
    "1111000100000101",
    "1111001000100101",
    "1111010001001100",
    "1111011011100101",
    "1111100101100000",
    "1111101101110001",
    "1111110101100011",
    "1111111111100010",
    "1111110001110000",
    "1111011101111101",
    "1111000111100010",
    "1110110011001111",
    "1110100110100100",
    "1110100101110100",
    "1110110010011101",
    "1111001010000111",
    "1111100111100111",
    "1111111011011000",
    "1111100100100000",
    "1111010111010101",
    "1111010101011111",
    "1111011110110101",
    "1111110001110101",
    "1111110100001100",
    "1111010110101101",
    "1110111001011011",
    "1110011111110000",
    "1110001100011001",
    "1110000001000010",
    "1101111101101110",
    "1110000000110000",
    "1110000111010011",
    "1110001110101000",
    "1110010100110011",
    "1110011001001011",
    "1110011100000010",
    "1110011110010110",
    "1110100001001101",
    "1110100101110110",
    "1110101101011110",
    "1110111001000110",
    "1111001001011101",
    "1111011110100110",
    "1111110111100111",
    "1111101101101001",
    "1111010100010111",
    "1110111111111011",
    "1110110011000000",
    "1110101110110011",
    "1110110010111001",
    "1110111101100011",
    "1111001100100000",
    "1111011101110101",
    "1111110000010010",
    "1111111100110111",
    "1111101010101000",
    "1111011010011000",
    "1111001101110111",
    "1111000110101111",
    "1111000101101010",
    "1111001010000110",
    "1111010010011101",
    "1111011100111000",
    "1111100111111111",
    "1111110011010110",
    "1111111111010011",
    "1111110011101100",
    "1111100101110110",
    "1111011000010110",
    "1111001101010001",
    "1111000111000011",
    "1111000111110001",
    "1111010000011100",
    "1111100000111001",
    "1111110111010110",
    "1111101111010110",
    "1111010111001001",
    "1111000011110011",
    "1110111000010001",
    "1110110110010110",
    "1110111110010111",
    "1111001111101110",
    "1111101001000001",
    "1111111000001001",
    "1111010111000001",
    "1110110111010101",
    "1110011100110010",
    "1110001010011000",
    "1110000001100100",
    "1110000001111101",
    "1110001001100111",
    "1110010110001001",
    "1110100101110111",
    "1110111000010000",
    "1111001101011001",
    "1111100101010010",
    "1111111110110110",
    "1111100111111111",
    "1111010010010100",
    "1111000010110110",
    "1110111011001110",
    "1110111011010011",
    "1111000001101001",
    "1111001100001111",
    "1111011001010011",
    "1111100111110010",
    "1111110111000111",
    "1111111001010000",
    "1111101010011100",
    "1111011101111101",
    "1111010101011011",
    "1111010001111110",
    "1111010011110100",
    "1111011010000001",
    "1111100010111011",
    "1111101100011110",
    "1111110100110110",
    "1111111010110100",
    "1111111101110110",
    "1111111110000100",
    "1111111011111101",
    "1111111000010100",
    "1111110011111111",
    "1111101111101100",
    "1111101100000010",
    "1111101001010010",
    "1111100111010111",
    "1111100101101001",
    "1111100010111001",
    "1111011101110011",
    "1111010101011101",
    "1111001010001100",
    "1110111101100001",
    "1110110001111000",
    "1110101001110010",
    "1110100111001011",
    "1110101010110111",
    "1110110100110110",
    "1111000100011101",
    "1111011000110100",
    "1111110000011100",
    "1111110110110100",
    "1111100000001000",
    "1111001110110110",
    "1111000101110001",
    "1111000110001101",
    "1111001111100100",
    "1111011111110001",
    "1111110100000010",
    "1111110110000101",
    "1111100000011010",
    "1111001100010110",
    "1110111011001110",
    "1110101110101110",
    "1110101000111100",
    "1110101011111000",
    "1110111000011101",
    "1111001101011001",
    "1111100111010101",
    "1111111110010101",
    "1111101000001000",
    "1111011000111001",
    "1111010001001101",
    "1111001111101110",
    "1111010001111011",
    "1111010101011111",
    "1111011000111110",
    "1111011100000101",
    "1111011111010010",
    "1111100011000101",
    "1111100111101110",
    "1111101101000001",
    "1111110010101011",
    "1111111000100001",
    "1111111110111010",
    "1111111001010000",
    "1111101111000011",
    "1111100001111000",
    "1111010010010000",
    "1111000001101011",
    "1110110010010010",
    "1110100101111110",
    "1110011101110011",
    "1110011001110010",
    "1110011001000110",
    "1110011010101010",
    "1110011101101001",
    "1110100001110001",
    "1110100111010011",
    "1110101110100011",
    "1110110111011111",
    "1111000001100001",
    "1111001011100101",
    "1111010100011000",
    "1111011010111100",
    "1111011110101011",
    "1111011111100100",
    "1111011110000000",
    "1111011010100010",
    "1111010101100111",
    "1111001111111000",
    "1111001010001110",
    "1111000101111110",
    "1111000100101110",
    "1111000111111001",
    "1111010000011100",
    "1111011110011100",
    "1111110001000010",
    "1111111001100110",
    "1111100100000001",
    "1111010000110110",
    "1111000010010010",
    "1110111001100000",
    "1110110110100111",
    "1110111000110101",
    "1110111111000111",
    "1111001000001110",
    "1111010011011010",
    "1111100000001100",
    "1111101110001110",
    "1111111101001101",
    "1111110011100111",
    "1111100101100000",
    "1111011001110010",
    "1111010001100110",
    "1111001101100110",
    "1111001101101011",
    "1111010001000010",
    "1111010110100000",
    "1111011101000000",
    "1111100011101100",
    "1111101010001101",
    "1111110000100100",
    "1111110110110011",
    "1111111100111010",
    "1111111101010101",
    "1111111000010111",
    "1111110100100000",
    "1111110001111011",
    "1111110000011011",
    "1111101111011100",
    "1111101110011010",
    "1111101100110100",
    "1111101010100111",
    "1111101000000010",
    "1111100101011011",
    "1111100010111110",
    "1111100000101100",
    "1111011110011011",
    "1111011100000101",
    "1111011001110101",
    "1111011000001001",
    "1111010111100011",
    "1111011000100101",
    "1111011011010100",
    "1111011111011110",
    "1111100100001110",
    "1111101000110101",
    "1111101100101001",
    "1111101111100011",
    "1111110010000100",
    "1111110101001000",
    "1111111010000000",
    "1111111110010000",
    "1111110011010111",
    "1111100110000001",
    "1111010111111110",
    "1111001011101010",
    "1111000011011100",
    "1111000000111011",
    "1111000100101001",
    "1111001110001101",
    "1111011100101011",
    "1111101110111101",
    "1111111100000000",
    "1111100101101110",
    "1111010000001000",
    "1110111101111011",
    "1110110001111001",
    "1110101110011001",
    "1110110100111011",
    "1111000101011010",
    "1111011101111111",
    "1111111011001101",
    "1111100111001111",
    "1111001101101011",
    "1110111011001001",
    "1110110001001111",
    "1110101111110110",
    "1110110101111011",
    "1111000001110110",
    "1111010010001111",
    "1111100101110111",
    "1111111011011001",
    "1111101111001000",
    "1111011100000111",
    "1111001101110111",
    "1111000101111011",
    "1111000100101001",
    "1111001000110000",
    "1111010000000000",
    "1111010111100101",
    "1111011101001001",
    "1111011111010110",
    "1111011110001010",
    "1111011010100110",
    "1111010110010010",
    "1111010010101100",
    "1111010001001101",
    "1111010011000110",
    "1111011001011000",
    "1111100100011010",
    "1111110011001101",
    "1111111100010110",
    "1111101101010100",
    "1111100010011100",
    "1111011101010010",
    "1111011101101101",
    "1111100001110110",
    "1111100110111111",
    "1111101010101110",
    "1111101100001110",
    "1111101100110001",
    "1111101110110110",
    "1111110100110100",
    "1111111111100000",
    "1111110010011110",
    "1111100100011101",
    "1111011010010100",
    "1111010111000100",
    "1111011011110000",
    "1111100111100000",
    "1111111000100010",
    "1111110011000010",
    "1111011101001010",
    "1111000111110001",
    "1110110101001000",
    "1110100111101111",
    "1110100001100110",
    "1110100011101110",
    "1110101101010110",
    "1110111011111100",
    "1111001100001100",
    "1111011011011001",
    "1111101001010000",
    "1111110111111101",
    "1111110101011011",
    "1111011101001010",
    "1111000000010111",
    "1110100011001000",
    "1110001010111000",
    "1101111100010011",
    "1101111001000111",
    "1101111111011001",
    "1110001010110010",
    "1110010110101000",
    "1110100000000101",
    "1110100110110111",
    "1110101100100001",
    "1110110011001011",
    "1110111100010111",
    "1111000111111010",
    "1111010100010010",
    "1111011111001010",
    "1111100110010010",
    "1111101000010110",
    "1111100101011111",
    "1111011110111011",
    "1111010110011111",
    "1111001101111011",
    "1111000111000011",
    "1111000011011111",
    "1111000100110011",
    "1111001011110111",
    "1111011000100011",
    "1111101001100111",
    "1111111100110011",
    "1111110000011101",
    "1111100000100001",
    "1111010100110100",
    "1111001101110010",
    "1111001010110101",
    "1111001010110111",
    "1111001100111000",
    "1111010000010100",
    "1111010101001011",
    "1111011011111000",
    "1111100101000001",
    "1111110001000011",
    "1111111111111011",
    "1111101111000101",
    "1111011101100011",
    "1111001101100001",
    "1111000001010000",
    "1110111010110101",
    "1110111011111000",
    "1111000101011111",
    "1111010111101100",
    "1111110001000010",
    "1111110001011111",
    "1111010100001011",
    "1110111011011001",
    "1110101010101011",
    "1110100011111000",
    "1110100110011101",
    "1110110000000000",
    "1110111101101110",
    "1111001110010111",
    "1111100010010100",
    "1111111010011010",
    "1111101001100001",
    "1111001100000010",
    "1110110001001100",
    "1110011101101000",
    "1110010100111001",
    "1110010111110111",
    "1110100100100000",
    "1110110111000001",
    "1111001011000100",
    "1111011101010010",
    "1111101011101010",
    "1111110101000101",
    "1111111000110011",
    "1111110110010001",
    "1111101101001011",
    "1111011110000100",
    "1111001010101000",
    "1110110101100111",
    "1110100010011100",
    "1110010100000101",
    "1110001100010111",
    "1110001011011011",
    "1110010000000010",
    "1110011000011010",
    "1110100010111011",
    "1110101110101101",
    "1110111011001111",
    "1111001000011110",
    "1111010110011111",
    "1111100101010101",
    "1111110101001101",
    "1111111001011100",
    "1111100110010110",
    "1111010001100110",
    "1110111100010011",
    "1110101000100000",
    "1110011001000111",
    "1110010000101011",
    "1110010000011100",
    "1110010111111110",
    "1110100100110011",
    "1110110011010111",
    "1111000000001101",
    "1111001000111111",
    "1111001101001010",
    "1111001101101001",
    "1111001101000101",
    "1111001111111000",
    "1111011010000111",
    "1111101101011001",
    "1111111000000110",
    "1111011011011101",
    "1111000010111110",
    "1110110100000110",
    "1110110001110011",
    "1110111011011000",
    "1111001101000111",
    "1111100010100100",
    "1111111000001101",
    "1111110011100100",
    "1111100001000010",
    "1111010000011001",
    "1111000010011001",
    "1110111000101101",
    "1110110101101111",
    "1110111011100001",
    "1111001010100000",
    "1111100000110011",
    "1111111010010110",
    "1111101101110101",
    "1111011011111101",
    "1111010010000101",
    "1111001111111111",
    "1111010011110011",
    "1111011011010100",
    "1111100100101010",
    "1111101110101000",
    "1111111000110111",
    "1111111100101000",
    "1111110010000110",
    "1111101000000000",
    "1111011111011010",
    "1111011001101010",
    "1111011000000100",
    "1111011011101011",
    "1111100100110001",
    "1111110010101001",
    "1111111100001100",
    "1111101001110101",
    "1111011000010001",
    "1111001001001001",
    "1110111101100110",
    "1110110110011111",
    "1110110100001000",
    "1110110110111001",
    "1110111111010010",
    "1111001110000010",
    "1111100011111001",
    "1111111111010000",
    "1111011101010100",
    "1110111001111001",
    "1110011001100111",
    "1110000000110110",
    "1101110010010111",
    "1101101110111010",
    "1101110101010000",
    "1110000010110110",
    "1110010101000101",
    "1110101010000010",
    "1111000000111011",
    "1111011001010101",
    "1111110010011101",
    "1111110101001011",
    "1111011111110001",
    "1111001111011100",
    "1111000101100000",
    "1111000010001010",
    "1111000100001011",
    "1111001001100011",
    "1111010000010101",
    "1111010111011101",
    "1111011111000111",
    "1111101000000100",
    "1111110011000001",
    "1111111111110000",
    "1111110011001011",
    "1111101000100111",
    "1111100011111001",
    "1111100111111100",
    "1111110101110000",
    "1111110100001100",
    "1111011001111111",
    "1111000000111101",
    "1110101110001101",
    "1110100101011010",
    "1110100111100111",
    "1110110011010010",
    "1111000101000110",
    "1111011001001001",
    "1111101100011101",
    "1111111110000010",
    "1111110001001101",
    "1111011111111101",
    "1111001101101101",
    "1110111011111010",
    "1110101101111010",
    "1110100111110100",
    "1110101100111000",
    "1110111101110010",
    "1111010111110100",
    "1111110101101110",
    "1111101110100001",
    "1111011001111010",
    "1111001110111011",
    "1111001101010111",
    "1111010010111110",
    "1111011100100000",
    "1111100110111111",
    "1111110000100001",
    "1111111000010001",
    "1111111110001101",
    "1111111101011111",
    "1111111010101111",
    "1111111001010000",
    "1111111000011001",
    "1111110110111010",
    "1111110011000100",
    "1111101010111110",
    "1111011101001010",
    "1111001001011101",
    "1110110001001101",
    "1110010111011010",
    "1101111111110000",
    "1101101101110000",
    "1101100011100010",
    "1101100001011001",
    "1101100101100010",
    "1101101101001001",
    "1101110101001001",
    "1101111011010100",
    "1101111110110101",
    "1110000000001101",
    "1110000001011111",
    "1110000110000000",
    "1110010000111101",
    "1110100011111000",
    "1110111101011100",
    "1111011001101101",
    "1111110011001111",
    "1111111010111010",
    "1111110011111110",
    "1111111000000100",
    "1111111011100100",
    "1111101011010101",
    "1111011011101011",
    "1111001111111011",
    "1111001001111001",
    "1111001010001111",
    "1111010000110101",
    "1111011100111000",
    "1111101101010001",
    "1111111111100101",
    "1111101100001011",
    "1111011011001001",
    "1111001111010010",
    "1111001010101101",
    "1111001110011011",
    "1111011001111111",
    "1111101011111011",
    "1111111101110011",
    "1111100101110001",
    "1111001110011110",
    "1110111010100000",
    "1110101011110010",
    "1110100011001111",
    "1110100000101110",
    "1110100011000110",
    "1110101000111100",
    "1110110000111001",
    "1110111010011101",
    "1111000101100101",
    "1111010010110011",
    "1111100010011100",
    "1111110100011011",
    "1111111000001001",
    "1111100100111110",
    "1111010100000110",
    "1111000111100101",
    "1111000001000101",
    "1111000001011100",
    "1111001000011110",
    "1111010101000101",
    "1111100101010011",
    "1111110110101000",
    "1111111001110000",
    "1111101110101101",
    "1111101010010101",
    "1111101101100100",
    "1111110111110010",
    "1111111000111001",
    "1111100111010100",
    "1111010110010010",
    "1111001000001000",
    "1110111110010111",
    "1110111001011101",
    "1110111000111100",
    "1110111011110111",
    "1111000001001000",
    "1111000111110111",
    "1111001111011110",
    "1111010111110010",
    "1111100001001000",
    "1111101100000100",
    "1111111001001100",
    "1111110111100100",
    "1111100111011000",
    "1111011000001110",
    "1111001100100011",
    "1111000110011111",
    "1111000111000011",
    "1111001110000100",
    "1111011001111111",
    "1111101000101110",
    "1111111000100001",
    "1111110111010101",
    "1111100110111000",
    "1111010101111100",
    "1111000101010011",
    "1110110110110111",
    "1110101101100001",
    "1110101100010100",
    "1110110101010011",
    "1111001000010110",
    "1111100010111110",
    "1111111111000000",
    "1111100010100010",
    "1111001011100101",
    "1110111100100101",
    "1110110110000011",
    "1110110111011011",
    "1110111111110000",
    "1111001110010001",
    "1111100010010101",
    "1111111010110110",
    "1111101010011000",
    "1111010000101110",
    "1110111100000010",
    "1110101111100100",
    "1110101100111100",
    "1110110011100001",
    "1111000000101110",
    "1111010000110011",
    "1111011111110101",
    "1111101010100110",
    "1111101111000010",
    "1111101100010000",
    "1111100010110001",
    "1111010100000110",
    "1111000010101110",
    "1110110001011110",
    "1110100011010011",
    "1110011010100110",
    "1110011000110111",
    "1110011110011111",
    "1110101010110000",
    "1110111100001010",
    "1111010000100111",
    "1111100101110010",
    "1111111001011011",
    "1111110110010101",
    "1111101010111101",
    "1111100101000000",
    "1111100100010000",
    "1111100111110110",
    "1111101110010100",
    "1111110110001001",
    "1111111101111010",
    "1111111011011111",
    "1111110111000100",
    "1111110101100000",
    "1111110111010101",
    "1111111100110000",
    "1111111010100101",
    "1111101111101101",
    "1111100011111100",
    "1111011000111001",
    "1111001111111111",
    "1111001010010100",
    "1111001000011000",
    "1111001001111101",
    "1111001110011001",
    "1111010100110001",
    "1111011100001110",
    "1111100100011000",
    "1111101110000101",
    "1111111011000110",
    "1111110010111001",
    "1111011011100110",
    "1111000000101011",
    "1110100101101010",
    "1110001111000111",
    "1110000001010010",
    "1101111110100011",
    "1110000110100101",
    "1110010110101010",
    "1110101010101000",
    "1110111110011001",
    "1111001110110110",
    "1111011010100010",
    "1111100001010101",
    "1111100100010011",
    "1111100100111001",
    "1111100100011101",
    "1111100011111000",
    "1111100011100010",
    "1111100011011111",
    "1111100011100010",
    "1111100011100010",
    "1111100011011010",
    "1111100011001000",
    "1111100010110110",
    "1111100010101111",
    "1111100011000001",
    "1111100011110100",
    "1111100100111011",
    "1111100110000011",
    "1111100110101110",
    "1111100110011111",
    "1111100101001000",
    "1111100010101001",
    "1111011111010100",
    "1111011011101011",
    "1111011000001100",
    "1111010101001001",
    "1111010010100010",
    "1111010000010001",
    "1111001110010010",
    "1111001100111101",
    "1111001100110010",
    "1111001110010110",
    "1111010001111001",
    "1111010111000001",
    "1111011100100101",
    "1111100001010000",
    "1111100100000110",
    "1111100100110011",
    "1111100011101110",
    "1111100001100110",
    "1111011111000100",
    "1111011100010110",
    "1111011001010000",
    "1111010101100000",
    "1111010000111011",
    "1111001011101111",
    "1111000110011000",
    "1111000001011001",
    "1110111100111010",
    "1110111000110101",
    "1110110100101111",
    "1110110000011001",
    "1110101011110101",
    "1110100111100011",
    "1110100100010101",
    "1110100010110110",
    "1110100011100100",
    "1110100110101010",
    "1110101100000100",
    "1110110011101001",
    "1110111101000000",
    "1111000111011111",
    "1111010001111101",
    "1111011010111111",
    "1111100001001010",
    "1111100011100010",
    "1111100010000011",
    "1111011101100100",
    "1111010111110111",
    "1111010011000001",
    "1111010001001010",
    "1111010011110110",
    "1111011011111101",
    "1111101001110001",
    "1111111100110100",
    "1111101100000001",
    "1111010010111001",
    "1110111010100010",
    "1110100101110001",
    "1110010111000011",
    "1110001111110110",
    "1110010000010010",
    "1110010111000110",
    "1110100001111110",
    "1110101110000000",
    "1110111000010000",
    "1110111110001111",
    "1110111110001111",
    "1110110111100111",
    "1110101011000110",
    "1110011010110000",
    "1110001001101101",
    "1101111011001010",
    "1101110001110000",
    "1101101110011110",
    "1101110000110101",
    "1101110110111111",
    "1101111110110101",
    "1110000111111110",
    "1110010100100010",
    "1110100111001101",
    "1111000001000011",
    "1111100000000010",
    "1111111111000110",
    "1111100111110011",
    "1111011001110101",
    "1111011001000010",
    "1111100011000110",
    "1111110010110010",
    "1111111101101010",
    "1111110010010111",
    "1111101011111110",
    "1111101000001011",
    "1111100011011010",
    "1111011010100010",
    "1111001100111000",
    "1110111100110011",
    "1110101110011100",
    "1110100110011010",
    "1110100111110101",
    "1110110011001010",
    "1111000101111011",
    "1111011100000100",
    "1111110001010011",
    "1111111101110111",
    "1111110011111001",
    "1111110001111000",
    "1111110111100000",
    "1111111100101101",
    "1111101101001011",
    "1111011100011100",
    "1111001100111101",
    "1111000000100110",
    "1110111000100011",
    "1110110101000110",
    "1110110101100010",
    "1110111000101010",
    "1110111101010001",
    "1111000010100010",
    "1111001000010000",
    "1111001110100011",
    "1111010101101110",
    "1111011101111000",
    "1111100110101010",
    "1111101111100000",
    "1111110111110010",
    "1111111111000001",
    "1111111011001001",
    "1111110111001110",
    "1111110101110100",
    "1111110111011100",
    "1111111100010101",
    "1111111011111110",
    "1111110010110100",
    "1111101001110110",
    "1111100010111001",
    "1111011111011100",
    "1111100000001101",
    "1111100100111110",
    "1111101100100001",
    "1111110101100011",
    "1111111110111011",
    "1111110111111011",
    "1111101111010001",
    "1111100111000101",
    "1111011111011001",
    "1111011000010110",
    "1111010010011111",
    "1111001110010111",
    "1111001100011001",
    "1111001100110000",
    "1111001111001100",
    "1111010011001101",
    "1111011000011101",
    "1111011111000111",
    "1111100111111000",
    "1111110011110111",
    "1111111100001100",
    "1111101000101100",
    "1111010011011111",
    "1110111111100100",
    "1110110000001101",
    "1110100111101010",
    "1110100110110010",
    "1110101100110111",
    "1110111000000110",
    "1111000110011000",
    "1111010101110010",
    "1111100100101111",
    "1111110001110100",
    "1111111011011110",
    "1111111111110101",
    "1111111110011100",
    "1111110101111111",
    "1111100111101011",
    "1111010101110111",
    "1111000011110110",
    "1110110100111001",
    "1110101011101011",
    "1110101001100010",
    "1110101110011001",
    "1110111001011000",
    "1111001001001011",
    "1111011100001111",
    "1111110000111010",
    "1111111010101001",
    "1111101000011000",
    "1111011001110010",
    "1111001111101110",
    "1111001010000001",
    "1111000111100101",
    "1111000110110110",
    "1111000110010000",
    "1111000100110011",
    "1111000010011001",
    "1110111111101001",
    "1110111101101110",
    "1110111101110101",
    "1111000000110101",
    "1111000111010000",
    "1111010001100001",
    "1111100000000111",
    "1111110011001000",
    "1111110110001000",
    "1111011101111010",
    "1111000111011000",
    "1110110110000100",
    "1110101100100001",
    "1110101011011000",
    "1110110001001111",
    "1110111011011000",
    "1111000111001001",
    "1111010011101010",
    "1111100001110100",
    "1111110011010001",
    "1111110111001001",
    "1111011110110011",
    "1111000111000011",
    "1110110100001110",
    "1110101010000001",
    "1110101001101111",
    "1110110010000010",
    "1110111111100110",
    "1111001110111111",
    "1111011101110011",
    "1111101011100011",
    "1111111000111000",
    "1111111001100001",
    "1111101100000110",
    "1111100000101001",
    "1111011001110100",
    "1111011001111111",
    "1111100010001101",
    "1111110001011101",
    "1111111011001010",
    "1111100111100010",
    "1111010111001101",
    "1111001100100101",
    "1111001000100011",
    "1111001010101111",
    "1111010001111011",
    "1111011100101000",
    "1111101001011110",
    "1111110111000111",
    "1111111011101110",
    "1111110000011010",
    "1111101000001010",
    "1111100011111100",
    "1111100100001011",
    "1111101000110001",
    "1111110001000110",
    "1111111100001110",
    "1111110110111011",
    "1111101001100111",
    "1111011100111111",
    "1111010001111110",
    "1111001001010001",
    "1111000011001101",
    "1110111111101011",
    "1110111110010110",
    "1110111110110101",
    "1111000000111110",
    "1111000101001110",
    "1111001100010111",
    "1111010111010000",
    "1111100110000110",
    "1111111000001111",
    "1111110100000001",
    "1111100001001010",
    "1111010001100100",
    "1111000111000100",
    "1111000010011001",
    "1111000011000001",
    "1111000111110010",
    "1111001111000111",
    "1111010111100111",
    "1111100000010001",
    "1111101000011011",
    "1111101111110101",
    "1111110110011011",
    "1111111100001001",
    "1111111111000000",
    "1111111011010011",
    "1111111001001010",
    "1111111001001010",
    "1111111100000100",
    "1111111101100001",
    "1111110011101001",
    "1111100111000111",
    "1111011001100010",
    "1111001100111010",
    "1111000011001101",
    "1110111101101110",
    "1110111100111000",
    "1111000000001000",
    "1111000110010110",
    "1111001110100001",
    "1111011000011101",
    "1111100100101110",
    "1111110100000010",
    "1111111001101101",
    "1111100110001110",
    "1111010100100100",
    "1111001000101010",
    "1111000110011010",
    "1111010000000101",
    "1111100101001101",
    "1111111101100101",
    "1111011101100110",
    "1111000000011001",
    "1110101010011101",
    "1110011110000000",
    "1110011010111100",
    "1110011111010100",
    "1110101000110100",
    "1110110110010000",
    "1111000111111010",
    "1111011110101011",
    "1111111010100110",
    "1111100110001000",
    "1111000111000100",
    "1110101100010110",
    "1110011001001001",
    "1110001110011111",
    "1110001011001111",
    "1110001100100110",
    "1110001111101001",
    "1110010010001111",
    "1110010011111000",
    "1110010101000110",
    "1110010110111110",
    "1110011010001100",
    "1110011111001100",
    "1110100110011101",
    "1110110001000000",
    "1111000000000111",
    "1111010100011101",
    "1111101101010110",
    "1111110111110110",
    "1111011111001111",
    "1111001101000100",
    "1111000100001000",
    "1111000100101001",
    "1111001100000100",
    "1111010110100000",
    "1111100000010101",
    "1111100111010111",
    "1111101011001001",
    "1111101100011111",
    "1111101100100111",
    "1111101100010110",
    "1111101011101101",
    "1111101010000111",
    "1111100111000110",
    "1111100010100100",
    "1111011101000111",
    "1111010111110001",
    "1111010011010111",
    "1111010000001111",
    "1111001110011001",
    "1111001101101110",
    "1111001110100001",
    "1111010001101011",
    "1111011000100010",
    "1111100100101001",
    "1111110110101011",
    "1111110001111000",
    "1111010111001101",
    "1110111100100110",
    "1110100101101110",
    "1110010101100101",
    "1110001101110011",
    "1110001110011001",
    "1110010110000100",
    "1110100010111001",
    "1110110010111001",
    "1111000100010111",
    "1111010101110010",
    "1111100101101010",
    "1111110010011010",
    "1111111010101111",
    "1111111101111010",
    "1111111100000011",
    "1111110110001100",
    "1111101101111110",
    "1111100101001000",
    "1111011101000111",
    "1111010110101100",
    "1111010001110011",
    "1111001101111011",
    "1111001010010100",
    "1111000110011111",
    "1111000010011001",
    "1110111110100001",
    "1110111011111101",
    "1110111011111000",
    "1110111111100100",
    "1111000111110010",
    "1111010100011100",
    "1111100100100100",
    "1111110110010011",
    "1111111000100011",
    "1111101010001010",
    "1111100000000010",
    "1111011010101101",
    "1111011001110000",
    "1111011100001100",
    "1111100000101100",
    "1111100101111110",
    "1111101010111111",
    "1111101110111011",
    "1111110001010101",
    "1111110001111010",
    "1111110000101001",
    "1111101101101110",
    "1111101001011110",
    "1111100100010011",
    "1111011110101001",
    "1111011000111100",
    "1111010011011010",
    "1111001110010100",
    "1111001001111010",
    "1111000110100101",
    "1111000100110110",
    "1111000101001101",
    "1111001000001110",
    "1111001110010100",
    "1111010111111110",
    "1111100101101110",
    "1111111000010010",
    "1111110000000001",
    "1111010011111110",
    "1110110101101110",
    "1110011000110010",
    "1110000001001100",
    "1101110010010101",
    "1101101101111101",
    "1101110011110100",
    "1110000010000000",
    "1110010101111110",
    "1110101101011011",
    "1111000110101101",
    "1111100000101001",
    "1111111001110000",
    "1111101111111101",
    "1111011111000010",
    "1111010110000100",
    "1111010111001000",
    "1111100010101011",
    "1111110110111100",
    "1111110000000000",
    "1111010111010001",
    "1111000011011111",
    "1110110111101100",
    "1110110100101110",
    "1110111001100000",
    "1111000011101111",
    "1111010000111110",
    "1111011111010100",
    "1111101101100011",
    "1111111010110110",
    "1111111001101001",
    "1111110001001111",
    "1111101101001110",
    "1111101110011101",
    "1111110100111111",
    "1111111111110001",
    "1111110011001000",
    "1111100110000110",
    "1111011011001100",
    "1111010011100111",
    "1111001111011110",
    "1111001110000000",
    "1111001110010001",
    "1111001111100001",
    "1111010001011010",
    "1111010011111011",
    "1111010111000110",
    "1111011010110100",
    "1111011110110101",
    "1111100010110110",
    "1111100110011110",
    "1111101001011111",
    "1111101011111010",
    "1111101101111001",
    "1111101111101100",
    "1111110001011100",
    "1111110011001010",
    "1111110100110110",
    "1111110110100000",
    "1111111000011010",
    "1111111011000000",
    "1111111110111111",
    "1111111011000100",
    "1111110010111100",
    "1111101000110101",
    "1111011101110010",
    "1111010011011000",
    "1111001011101010",
    "1111001000011000",
    "1111001010110111",
    "1111010011100100",
    "1111100001101110",
    "1111110011011101",
    "1111111001111001",
    "1111101001001100",
    "1111011100101101",
    "1111010101110100",
    "1111010100100000",
    "1111010111100101",
    "1111011101000100",
    "1111100010111011",
    "1111100111110010",
    "1111101011001001",
    "1111101101011100",
    "1111101111101011",
    "1111110010110111",
    "1111110111101011",
    "1111111110001011",
    "1111111010000010",
    "1111110001110101",
    "1111101010000010",
    "1111100011010111",
    "1111011110010110",
    "1111011011010011",
    "1111011010011001",
    "1111011011101010",
    "1111011110111000",
    "1111100011100010",
    "1111101000110011",
    "1111101101100101",
    "1111110000101100",
    "1111110001001001",
    "1111101110011111",
    "1111101000111110",
    "1111100001011001",
    "1111011001000111",
    "1111010001101001",
    "1111001100010100",
    "1111001010000010",
    "1111001011000110",
    "1111001111000111",
    "1111010101001101",
    "1111011100010110",
    "1111100011010000",
    "1111101000111011",
    "1111101100011111",
    "1111101101011110",
    "1111101011101111",
    "1111100111010001",
    "1111100000001101",
    "1111010110100010",
    "1111001010000010",
    "1110111010011000",
    "1110100111100011",
    "1110010010010101",
    "1101111100001111",
    "1101100111100111",
    "1101010110111110",
    "1101001100010110",
    "1101001000110010",
    "1101001011110111",
    "1101010011110001",
    "1101011110001010",
    "1101101000101100",
    "1101110001101011",
    "1101111000011011",
    "1101111101010001",
    "1110000001000101",
    "1110000101001000",
    "1110001010011110",
    "1110010001011111",
    "1110011001100000",
    "1110100001000010",
    "1110100110010011",
    "1110101000010011",
    "1110100111000001",
    "1110100011101110",
    "1110100000111101",
    "1110100001101100",
    "1110101000101100",
    "1110110111011011",
    "1111001101101001",
    "1111101001000101",
    "1111111010000010",
    "1111100000001101",
    "1111001101010001",
    "1111000011011101",
    "1111000010110110",
    "1111001001100010",
    "1111010100100101",
    "1111100001000101",
    "1111101100101110",
    "1111110110010010",
    "1111111101001110",
    "1111111110100001",
    "1111111100111001",
    "1111111101101011",
    "1111111111011100",
    "1111111011001111",
    "1111110110111000",
    "1111110100000100",
    "1111110100110011",
    "1111111010110110",
    "1111111000110101",
    "1111100111000010",
    "1111010010001000",
    "1110111101101000",
    "1110101101000111",
    "1110100011001101",
    "1110100000110001",
    "1110100100110111",
    "1110101101001100",
    "1110110111010001",
    "1111000001110110",
    "1111001101011001",
    "1111011011100011",
    "1111101101110100",
    "1111111011110111",
    "1111100011101100",
    "1111001101001111",
    "1110111100001010",
    "1110110010111011",
    "1110110001101100",
    "1110110111000001",
    "1111000000110110",
    "1111001101110010",
    "1111011101101101",
    "1111110001000001",
    "1111111000100111",
    "1111100001000101",
    "1111001011101000",
    "1110111011111101",
    "1110110100111100",
    "1110110111101101",
    "1111000011010010",
    "1111010101000110",
    "1111101001111100",
    "1111111111001000",
    "1111101101001011",
    "1111011100001110",
    "1111001110101110",
    "1111000101100111",
    "1111000001100110",
    "1111000010110110",
    "1111001000101100",
    "1111010001011100",
    "1111011010110100",
    "1111100010100110",
    "1111100111010100",
    "1111101000101101",
    "1111100111100010",
    "1111100101000001",
    "1111100010001010",
    "1111011111001100",
    "1111011011110000",
    "1111010111000100",
    "1111010000100110",
    "1111001000010110",
    "1110111111010001",
    "1110110110110110",
    "1110110000111101",
    "1110101111010010",
    "1110110011000101",
    "1110111100110010",
    "1111001011111111",
    "1111011111101001",
    "1111110101111010",
    "1111110011011101",
    "1111011110110110",
    "1111001110001111",
    "1111000010111001",
    "1110111101010100",
    "1110111101010001",
    "1111000001111001",
    "1111001010001100",
    "1111010101001101",
    "1111100010010100",
    "1111110001001000",
    "1111111110011101",
    "1111101100101101",
    "1111011010010001",
    "1111001000010101",
    "1110111000100011",
    "1110101100101011",
    "1110100101110111",
    "1110100100100111",
    "1110101000011010",
    "1110101111111101",
    "1110111001110010",
    "1111000100100100",
    "1111001111010100",
    "1111011001010110",
    "1111100001111000",
    "1111100111111111",
    "1111101010011101",
    "1111101000001111",
    "1111100000100110",
    "1111010011101111",
    "1111000011000001",
    "1110110000110101",
    "1110100000000011",
    "1110010011100100",
    "1110001101011001",
    "1110001110100100",
    "1110010111000110",
    "1110100110010000",
    "1110111010110010",
    "1111010010110001",
    "1111101011101011",
    "1111111101010110",
    "1111101011010010",
    "1111100000010010",
    "1111011101011100",
    "1111100010100110",
    "1111101110011011",
    "1111111111001000",
    "1111101101000001",
    "1111010111101100",
    "1111000010001101",
    "1110101110001001",
    "1110011101000111",
    "1110010000101011",
    "1110001001101111",
    "1110001000011011",
    "1110001011110010",
    "1110010001111101",
    "1110011000101101",
    "1110011110001101",
    "1110100001100100",
    "1110100010110100",
    "1110100011000011",
    "1110100011100100",
    "1110100101110110",
    "1110101011001100",
    "1110110100110100",
    "1111000011101001",
    "1111010111101111",
    "1111101111111001",
    "1111110110010111",
    "1111011110011110",
    "1111001011100101",
    "1110111111110000",
    "1110111011010001",
    "1110111100011100",
    "1111000000011110",
    "1111000100011101",
    "1111000110100100",
    "1111000110101100",
    "1111000111000011",
    "1111001011001111",
    "1111010110100101",
    "1111101010001101",
    "1111111011110000",
    "1111011111111011",
    "1111000111111010",
    "1110111000101101",
    "1110110100111100",
    "1110111100010100",
    "1111001100001100",
    "1111100000110011",
    "1111110110010110",
    "1111110110001111",
    "1111100111011011",
    "1111011110111010",
    "1111011101111101",
    "1111100101010101",
    "1111110100110010",
    "1111110101011001",
    "1111011100011011",
    "1111000100001000",
    "1110110000011111",
    "1110100100001101",
    "1110100000000101",
    "1110100010110011",
    "1110101001101010",
    "1110110001110011",
    "1110111000111100",
    "1110111101111000",
    "1111000000011001",
    "1111000001001010",
    "1111000001101001",
    "1111000011101110",
    "1111001000110111",
    "1111010001100100",
    "1111011100110000",
    "1111100111111110",
    "1111110000001010",
    "1111110010100000",
    "1111101101011001",
    "1111100001000011",
    "1111001111011110",
    "1110111011110000",
    "1110101001011001",
    "1110011011001110",
    "1110010011001011",
    "1110010010010000",
    "1110011000101010",
    "1110100110011101",
    "1110111011100000",
    "1111010111000110",
    "1111110111011011",
    "1111100110100000",
    "1111000110100111",
    "1110101100011100",
    "1110011010011000",
    "1110010000110110",
    "1110001110011100",
    "1110010000100110",
    "1110010100100111",
    "1110011000011101",
    "1110011011000110",
    "1110011100101101",
    "1110011110000010",
    "1110100000000101",
    "1110100011100010",
    "1110101000100000",
    "1110101110011001",
    "1110110100000110",
    "1110111000010001",
    "1110111001101010",
    "1110110111010110",
    "1110110001001100",
    "1110100111110010",
    "1110011100100110",
    "1110010001101110",
    "1110001001100011",
    "1110000110011010",
    "1110001010010011",
    "1110010110100101",
    "1110101011110101",
    "1111001001001011",
    "1111101011110111",
    "1111110000011011",
    "1111010000111000",
    "1110111010000111",
    "1110101110111101",
    "1110101111101110",
    "1110111010000110",
    "1111001010000010",
    "1111011011000111",
    "1111101001111010",
    "1111110101000110",
    "1111111101100111",
    "1111111010001001",
    "1111101111111001",
    "1111100010011111",
    "1111010010101111",
    "1111000011001010",
    "1110110111000001",
    "1110110001000011",
    "1110110010001101",
    "1110111001010110",
    "1111000011110100",
    "1111001110010111",
    "1111010110001110",
    "1111011001110101",
    "1111011001000001",
    "1111010100110111",
    "1111001111001000",
    "1111001001011110",
    "1111000101000000",
    "1111000010001111",
    "1111000001010010",
    "1111000010010000",
    "1111000101001110",
    "1111001010001100",
    "1111010000111000",
    "1111011000011011",
    "1111011111101000",
    "1111100101000001",
    "1111100111011110",
    "1111100110010011",
    "1111100001110011",
    "1111011011000111",
    "1111010100000001",
    "1111001110101001",
    "1111001100111000",
    "1111010000000010",
    "1111011000100010",
    "1111100101110001",
    "1111110110001010",
    "1111111000011100",
    "1111101000100010",
    "1111011100000111",
    "1111010100011100",
    "1111010001101011",
    "1111010010111110",
    "1111010111000001",
    "1111011100011011",
    "1111100010010101",
    "1111101000011111",
    "1111101111001001",
    "1111110110101110",
    "1111111111010101",
    "1111110111011010",
    "1111101110110010",
    "1111101000011100",
    "1111100110001011",
    "1111101001011110",
    "1111110010110001",
    "1111111110100100",
    "1111101100011100",
    "1111011001010110",
    "1111000111111010",
    "1110111010010110",
    "1110110010001000",
    "1110101111111011",
    "1110110011110110",
    "1110111101100110",
    "1111001100111100",
    "1111100001010000",
    "1111111001011111",
    "1111101100011101",
    "1111010011011101",
    "1110111110101001",
    "1110110000101100",
    "1110101011001100",
    "1110101110010010",
    "1110111000110111",
    "1111001001000001",
    "1111011100100101",
    "1111110001011101",
    "1111111010001111",
    "1111101000001110",
    "1111011001111010",
    "1111010000010010",
    "1111001011101101",
    "1111001011111101",
    "1111010000010111",
    "1111011000000100",
    "1111100010010000",
    "1111101110010001",
    "1111111011001100",
    "1111111000000101",
    "1111101101010001",
    "1111100110010101",
    "1111100101000011",
    "1111101010010111",
    "1111110101110011",
    "1111111010011011",
    "1111101001000100",
    "1111011000110010",
    "1111001011100101",
    "1111000010100010",
    "1110111101110101",
    "1110111101001110",
    "1111000000010101",
    "1111000111000011",
    "1111010001010000",
    "1111011110101110",
    "1111101111000000",
    "1111111110101001",
    "1111101011010000",
    "1111010111110101",
    "1111000101100010",
    "1110110101011011",
    "1110101000011110",
    "1110011111011001",
    "1110011010101010",
    "1110011010011011",
    "1110011110010111",
    "1110100101110111",
    "1110110000000111",
    "1110111100010110",
    "1111001010000111",
    "1111011001001011",
    "1111101001001110",
    "1111111001101001",
    "1111110110101010",
    "1111101001011100",
    "1111100000011110",
    "1111011101010100",
    "1111100000110011",
    "1111101010101100",
    "1111111001100011",
    "1111110100111010",
    "1111100011101010",
    "1111010101100101",
    "1111001101000101",
    "1111001011111101",
    "1111010011000001",
    "1111100001111000",
    "1111110110101010",
    "1111110001101111",
    "1111011011000111",
    "1111001000111001",
    "1110111101011001",
    "1110111001010001",
    "1110111011011110",
    "1111000001101100",
    "1111001001011011",
    "1111010000101011",
    "1111010110100100",
    "1111011010111101",
    "1111011110010100",
    "1111100001000011",
    "1111100011011010",
    "1111100101011000",
    "1111100110111010",
    "1111101000010000",
    "1111101010000110",
    "1111101101100000",
    "1111110011100101",
    "1111111101000100",
    "1111110110001010",
    "1111100111010111",
    "1111011000011101",
    "1111001011100110",
    "1111000010011100",
    "1110111101101001",
    "1110111100111100",
    "1110111111000111",
    "1111000010110100",
    "1111000111000011",
    "1111001011011001",
    "1111010000001010",
    "1111010101111001",
    "1111011101000010",
    "1111100101011111",
    "1111101110100110",
    "1111110111001000",
    "1111111101101100",
    "1111111110111111",
    "1111111111111101",
    "1111111010001111",
    "1111101111110011",
    "1111100001100010",
    "1111010001001000",
    "1111000000110110",
    "1110110011001011",
    "1110101010001100",
    "1110100111010000",
    "1110101010011110",
    "1110110011000101",
    "1110111111110000",
    "1111001111000000",
    "1111011111100110",
    "1111110000100110",
    "1111111110101011",
    "1111101111000110",
    "1111100001100100",
    "1111010111001001",
    "1111010000101011",
    "1111001110100001",
    "1111010000001101",
    "1111010100100111",
    "1111011001111101",
    "1111011110100100",
    "1111100001010101",
    "1111100001111110",
    "1111100001001010",
    "1111100000000101",
    "1111100000000010",
    "1111100001111110",
    "1111100110010011",
    "1111101100111010",
    "1111110101001000",
    "1111111110001010",
    "1111111000111000",
    "1111110000110011",
    "1111101010000111",
    "1111100100111011",
    "1111100001000000",
    "1111011101110010",
    "1111011010011011",
    "1111010110001110",
    "1111010000111110",
    "1111001010111111",
    "1111000101011000",
    "1111000001101100",
    "1111000001011010",
    "1111000101101010",
    "1111001110101110",
    "1111011011110101",
    "1111101011100001",
    "1111111011101101",
    "1111110101110011",
    "1111101010111100",
    "1111100100110110",
    "1111100011101100",
    "1111100110101010",
    "1111101100001000",
    "1111110010000111",
    "1111110110110101",
    "1111111001000111",
    "1111111000100111",
    "1111110101110101",
    "1111110001110101",
    "1111101101111101",
    "1111101011011100",
    "1111101011000010",
    "1111101100111000",
    "1111110000010110",
    "1111110100010111",
    "1111110111101001",
    "1111111001000100",
    "1111110111111110",
    "1111110100001010",
    "1111101101111011",
    "1111100101110100",
    "1111011100100110",
    "1111010011001011",
    "1111001010110000",
    "1111000100110110",
    "1111000010111101",
    "1111000110010110",
    "1111001111011010",
    "1111011101010100",
    "1111101101111011",
    "1111111110011000",
    "1111110100001110",
    "1111101100000110",
    "1111101010001000",
    "1111101101111111",
    "1111110110101011",
    "1111111100111001",
    "1111101101100101",
    "1111011011111000",
    "1111001000011000",
    "1110110100011010",
    "1110100001111101",
    "1110010011010111",
    "1110001010100110",
    "1110001000100000",
    "1110001100011001",
    "1110010100010010",
    "1110011101100001",
    "1110100101110001",
    "1110101011101101",
    "1110101111001100",
    "1110110001000101",
    "1110110010100111",
    "1110110100111011",
    "1110111000110100",
    "1110111110110011",
    "1111000111001001",
    "1111010010001000",
    "1111011111110000",
    "1111101111100011",
    "1111111111101101",
    "1111110000001100",
    "1111100100000110",
    "1111011101001110",
    "1111011011111111",
    "1111011111100011",
    "1111100110001000",
    "1111101101111011",
    "1111110101110000",
    "1111111101100011",
    "1111111001110000",
    "1111101110111101",
    "1111100001010010",
    "1111010001001010",
    "1111000000010100",
    "1110110001010101",
    "1110100110101101",
    "1110100001111110",
    "1110100011010000",
    "1110101001101000",
    "1110110011100010",
    "1110111111101001",
    "1111001101011011",
    "1111011100111010",
    "1111101110001010",
    "1111111111011110",
    "1111101101110101",
    "1111011111010001",
    "1111010110000001",
    "1111010011011111",
    "1111010111100111",
    "1111100001000111",
    "1111101101110000",
    "1111111011010110",
    "1111110111110111",
    "1111101101000100",
    "1111100100101111",
    "1111011111001101",
    "1111011100101010",
    "1111011101000100",
    "1111100000000011",
    "1111100100110001",
    "1111101010000000",
    "1111101110100100",
    "1111110001101001",
    "1111110011000011",
    "1111110011001010",
    "1111110010100101",
    "1111110001110101",
    "1111110000111111",
    "1111101111101100",
    "1111101101100000",
    "1111101010000100",
    "1111100101100010",
    "1111100000100011",
    "1111011100000111",
    "1111011001011101",
    "1111011001101011",
    "1111011101101101",
    "1111100101111001",
    "1111110010001000",
    "1111111110010011",
    "1111101100101100",
    "1111011010100010",
    "1111001001011011",
    "1110111010110000",
    "1110101111011111",
    "1110101000000110",
    "1110100100100101",
    "1110100100101001",
    "1110100111101111",
    "1110101101010110",
    "1110110101000110",
    "1110111111000000",
    "1111001011011001",
    "1111011010100000",
    "1111101011111000",
    "1111111110010000",
    "1111110000001011",
    "1111100001011111",
    "1111010110111111",
    "1111010001000011",
    "1111001110111000",
    "1111001110111000",
    "1111001111010111",
    "1111001111011111",
    "1111001111100011",
    "1111010000110001",
    "1111010100100000",
    "1111011011010001",
    "1111100100001000",
    "1111101100110111",
    "1111110010100011",
    "1111110010110110",
    "1111101100111011",
    "1111100001110110",
    "1111010100010101",
    "1111000111110001",
    "1110111111000010",
    "1110111011110111",
    "1110111110101001",
    "1111000110111001",
    "1111010011111100",
    "1111100101010101",
    "1111111010110110",
    "1111101100000000",
    "1111010000111001",
    "1110110110100111",
    "1110100000110001",
    "1110010010100110",
    "1110001101111101",
    "1110010010101100",
    "1110011110111111",
    "1110110000000011",
    "1111000011010111",
    "1111010111001110",
    "1111101010110110",
    "1111111101111110",
    "1111101111110000",
    "1111011111001101",
    "1111010001100001",
    "1111000111101101",
    "1111000010011101",
    "1111000001011111",
    "1111000011111000",
    "1111001000011010",
    "1111001101111111",
    "1111010100000011",
    "1111011010100011",
    "1111100001101011",
    "1111101001011111",
    "1111110001111001",
    "1111111010101001",
    "1111111100001110",
    "1111110010101011",
    "1111101000100111",
    "1111011110011110",
    "1111010101001110",
    "1111001110010010",
    "1111001011000010",
    "1111001100010111",
    "1111010010001000",
    "1111011011001001",
    "1111100101100101",
    "1111101111011100",
    "1111110111010100",
    "1111111100101001",
    "1111111111100111",
    "1111111111000001",
    "1111111110100111",
    "1111111110101101",
    "1111111111010000",
    "1111111111100010",
    "1111111101011011",
    "1111111010000000",
    "1111110100101010",
    "1111101100101100",
    "1111100001100110",
    "1111010011010101",
    "1111000010111000",
    "1110110010001011",
    "1110100011100111",
    "1110011001010101",
    "1110010100010011",
    "1110010100010111",
    "1110010111110111",
    "1110011100100001",
    "1110011111110101",
    "1110011111111010",
    "1110011011110000",
    "1110010011101001",
    "1110001000111001",
    "1101111101100001",
    "1101110011100111",
    "1101101100101011",
    "1101101001011000",
    "1101101001011101",
    "1101101011110111",
    "1101101111010110",
    "1101110010110001",
    "1101110101100101",
    "1101110111111010",
    "1101111010011011",
    "1101111110011111",
    "1110000110110111",
    "1110010110101100",
    "1110101111100100",
    "1111010000100110",
    "1111110101111101",
    "1111100110000001",
    "1111001001001001",
    "1110110111110001",
    "1110110011010010",
    "1110111001111100",
    "1111001000010101",
    "1111011010101101",
    "1111101110001000",
    "1111111111001001",
    "1111101110011000",
    "1111100000100110",
    "1111010110110010",
    "1111010010001000",
    "1111010011100110",
    "1111011011000100",
    "1111100111010110",
    "1111110110001000",
    "1111111011011011",
    "1111101111110010",
    "1111101000001101",
    "1111100100101010",
    "1111100100010101",
    "1111100110010011",
    "1111101010000100",
    "1111101111100011",
    "1111110111011000",
    "1111111101011011",
    "1111101110000011",
    "1111011010100101",
    "1111000100011111",
    "1110101110101101",
    "1110011100100110",
    "1110010001001000",
    "1110001110000100",
    "1110010011001111",
    "1110011111000000",
    "1110101110110101",
    "1111000001010100",
    "1111010111000001",
    "1111110001101101",
    "1111101101110111",
    "1111001001100010",
    "1110100101100101",
    "1110000111101111",
    "1101110101010101",
    "1101110001010100",
    "1101111010111100",
    "1110001110001010",
    "1110100101100111",
    "1110111100101011",
    "1111010000111011",
    "1111100001111101",
    "1111101111111110",
    "1111111010101110",
    "1111111110111000",
    "1111111110101000",
    "1111111010001000",
    "1111101011011111",
    "1111010111001101",
    "1111000000100100",
    "1110101011011011",
    "1110011010110000",
    "1110001111110011",
    "1110001010100000",
    "1110001010010001",
    "1110001110110011",
    "1110011000000110",
    "1110100110000110",
    "1110111000001001",
    "1111001100100110",
    "1111100001001101",
    "1111110011011010",
    "1111111110101011",
    "1111110101110110",
    "1111110001010101",
    "1111101111101000",
    "1111101111001010",
    "1111101110110100",
    "1111101110000111",
    "1111101100111001",
    "1111101011001111",
    "1111101001000101",
    "1111100110001110",
    "1111100010010100",
    "1111011101010110",
    "1111010111101100",
    "1111010010000010",
    "1111001100110010",
    "1111001000000001",
    "1111000011010010",
    "1110111110000101",
    "1110111000011000",
    "1110110010100111",
    "1110101101101110",
    "1110101010110101",
    "1110101010101101",
    "1110101101100001",
    "1110110010100110",
    "1110111000101010",
    "1110111110010111",
    "1111000010110011",
    "1111000101110111",
    "1111001000001011",
    "1111001010111100",
    "1111001111101000",
    "1111010111101010",
    "1111100100001010",
    "1111110101101010",
    "1111110011111110",
    "1111011010001001",
    "1110111111001010",
    "1110100101111001",
    "1110010001001000",
    "1110000010101100",
    "1101111011001110",
    "1101111001111111",
    "1101111101100100",
    "1110000100011100",
    "1110001101101101",
    "1110011001001110",
    "1110100111001110",
    "1110110111101101",
    "1111001001111010",
    "1111011100010001",
    "1111101100101011",
    "1111111001000110",
    "1111111111110000",
    "1111111110010011",
    "1111111110001101",
    "1111110111010110",
    "1111101110101110",
    "1111100101111110",
    "1111011110011110",
    "1111011001011001",
    "1111010111101101",
    "1111011001111101",
    "1111100000001000",
    "1111101001100101",
    "1111110101000000",
    "1111111111000010",
    "1111110100000101",
    "1111101011000111",
    "1111100100100010",
    "1111100000011001",
    "1111011110011100",
    "1111011110110001",
    "1111100001110100",
    "1111101000001011",
    "1111110010001010",
    "1111111111011110",
    "1111110001000000",
    "1111100000111101",
    "1111010010000101",
    "1111000101110001",
    "1110111100101110",
    "1110110111001101",
    "1110110101001001",
    "1110110110100101",
    "1110111011101011",
    "1111000100011101",
    "1111010000110101",
    "1111100000000000",
    "1111110000101101",
    "1111111110101110",
    "1111110000000110",
    "1111100100110100",
    "1111011101101011",
    "1111011010111000",
    "1111011100010100",
    "1111100001101110",
    "1111101010111100",
    "1111110111111111",
    "1111110111000011",
    "1111100010101110",
    "1111001100001111",
    "1110110101111110",
    "1110100010110100",
    "1110010101101010",
    "1110010000100110",
    "1110010100100010",
    "1110100001000101",
    "1110110100100000",
    "1111001100001100",
    "1111100100110110",
    "1111111011000100",
    "1111110100000111",
    "1111101011001001",
    "1111101011101100",
    "1111110110011100",
    "1111110101011010",
    "1111011010100000",
    "1110111100111000",
    "1110100001001000",
    "1110001011011001",
    "1101111110011011",
    "1101111010111111",
    "1101111111100110",
    "1110001001011000",
    "1110010101001101",
    "1110100000101001",
    "1110101010011001",
    "1110110010011100",
    "1110111001101010",
    "1111000001001111",
    "1111001010000110",
    "1111010100010000",
    "1111011111000010",
    "1111101001001101",
    "1111110001100110",
    "1111110111011001",
    "1111111010100100",
    "1111111011011110",
    "1111111010101110",
    "1111111000110110",
    "1111110110001100",
    "1111110010111011",
    "1111101111000011",
    "1111101010011111",
    "1111100101001101",
    "1111011111010100",
    "1111011001001011",
    "1111010011010011",
    "1111001110011001",
    "1111001010111100",
    "1111001001010011",
    "1111001001011101",
    "1111001011001001",
    "1111001110000000",
    "1111010001110011",
    "1111010110100101",
    "1111011100101110",
    "1111100101001011",
    "1111110001000111",
    "1111111110100011",
    "1111101010000011",
    "1111010010111011",
    "1110111011110111",
    "1110100111111110",
    "1110011001110111",
    "1110010010111110",
    "1110010011001000",
    "1110011000100011",
    "1110100000110110",
    "1110101001111010",
    "1110110010111110",
    "1110111100101011",
    "1111001000000011",
    "1111010101100101",
    "1111100100011111",
    "1111110010101011",
    "1111111101011100",
    "1111111101011100",
    "1111111110111010",
    "1111111010001101",
    "1111110000101000",
    "1111100111100010",
    "1111100001100010",
    "1111100000001101",
    "1111100011101110",
    "1111101011010100",
    "1111110101100101",
    "1111111111000010",
    "1111110011110100",
    "1111101001100000",
    "1111100000011001",
    "1111011000101000",
    "1111010010010111",
    "1111001101110010",
    "1111001011010110",
    "1111001011101000",
    "1111001111100110",
    "1111011000010001",
    "1111100110011111",
    "1111111010001111",
    "1111101101100111",
    "1111010011011100",
    "1110111010001111",
    "1110100101010111",
    "1110010111010101",
    "1110010001100110",
    "1110010100000000",
    "1110011100111111",
    "1110101010000100",
    "1110111000010110",
    "1111000101001101",
    "1111001110111000",
    "1111010100101001",
    "1111010110110111",
    "1111010110011111",
    "1111010100110001",
    "1111010010101111",
    "1111010001001111",
    "1111010000101011",
    "1111010001001100",
    "1111010010011101",
    "1111010100000000",
    "1111010101000101",
    "1111010101001001",
    "1111010011111011",
    "1111010001100111",
    "1111001111000101",
    "1111001101100110",
    "1111001110101011",
    "1111010011100111",
    "1111011100111111",
    "1111101010011001",
    "1111111010011001",
    "1111110101010001",
    "1111100111000111",
    "1111011101001010",
    "1111011000100011",
    "1111011001011000",
    "1111011111000000",
    "1111101000100100",
    "1111110101010110",
    "1111111010111010",
    "1111101000100011",
    "1111010100011101",
    "1111000000100100",
    "1110101111110000",
    "1110100101001000",
    "1110100011000000",
    "1110101010011000",
    "1110111010011101",
    "1111010000111110",
    "1111101011000001",
    "1111111010100101",
    "1111100010110011",
    "1111001111110110",
    "1111000011010011",
    "1110111101101110",
    "1110111110110011",
    "1111000101001011",
    "1111001110111011",
    "1111011001110100",
    "1111100011101111",
    "1111101011011101",
    "1111110000011101",
    "1111110011000111",
    "1111110100010000",
    "1111110100111111",
    "1111110110001101",
    "1111111000100100",
    "1111111100100111",
    "1111111100111100",
    "1111110011011000",
    "1111100110000011",
    "1111010100111100",
    "1111000001010111",
    "1110101101101000",
    "1110011100100001",
    "1110010000011010",
    "1110001010101000",
    "1110001011000010",
    "1110010000101011",
    "1110011010010001",
    "1110100111001110",
    "1110110111100011",
    "1111001011100011",
    "1111100010101110",
    "1111111011010001",
    "1111101101110001",
    "1111011011101111",
    "1111010000111001",
    "1111001110000111",
    "1111010010011010",
    "1111011011111101",
    "1111101001001100",
    "1111111001010111",
    "1111110011110001",
    "1111011111000010",
    "1111001010000100",
    "1110110111011101",
    "1110101001111010",
    "1110100011010111",
    "1110100100001000",
    "1110101010111100",
    "1110110101101001",
    "1111000010010100",
    "1111001111110000",
    "1111011101100110",
    "1111101011100011",
    "1111111000101111",
    "1111111100011001",
    "1111110110000011",
    "1111110101111110",
    "1111111100101100",
    "1111110110110100",
    "1111100111001110",
    "1111010111101101",
    "1111001011001110",
    "1111000011101100",
    "1111000001111101",
    "1111000110000110",
    "1111001111111111",
    "1111011111010010",
    "1111110011001111",
    "1111110101100100",
    "1111011101010111",
    "1111000110100101",
    "1110110011100001",
    "1110100101100100",
    "1110011101000111",
    "1110011001100101",
    "1110011001111100",
    "1110011101010111",
    "1110100011100111",
    "1110101100111000",
    "1110111001011000",
    "1111001000101111",
    "1111011001111001",
    "1111101011000101",
    "1111111010010010",
    "1111111010000011",
    "1111110010101100",
    "1111101111010001",
    "1111101110100100",
    "1111101110111110",
    "1111101111000110",
    "1111101110000000",
    "1111101011011000",
    "1111100111011111",
    "1111100010110100",
    "1111011101111111",
    "1111011001011000",
    "1111010100111100",
    "1111010000010101",
    "1111001011000010",
    "1111000100101111",
    "1110111101100001",
    "1110110101111110",
    "1110101111001101",
    "1110101010110000",
    "1110101001111111",
    "1110101101100110",
    "1110110101010101",
    "1111000000000011",
    "1111001100000001",
    "1111010111010001",
    "1111100000110101",
    "1111101001111001",
    "1111110101101101",
    "1111111000101100",
    "1111100000100100",
    "1111000100100000",
    "1110101001100111",
    "1110010101100000",
    "1110001100101110",
    "1110010000100011",
    "1110011110110000",
    "1110110011001101",
    "1111001001101101",
    "1111011111011110",
    "1111110011011000",
    "1111111011000010",
    "1111101100100100",
    "1111100010011001",
    "1111011110001100",
    "1111100001010010",
    "1111101011101000",
    "1111111011101101",
    "1111110001001100",
    "1111011110010010",
    "1111001110000010",
    "1111000001011111",
    "1110111000011010",
    "1110110001110011",
    "1110101100111101",
    "1110101001100101",
    "1110100111100111",
    "1110100110111111",
    "1110100111100000",
    "1110101001000100",
    "1110101011110101",
    "1110110000100111",
    "1110111000110100",
    "1111000110001000",
    "1111011001101011",
    "1111110011000110",
    "1111110000000101",
    "1111010011111000",
    "1110111100100000",
    "1110101101001111",
    "1110100111010001",
    "1110101001010011",
    "1110110000010001",
    "1110111000100101",
    "1110111111100001",
    "1111000011111000",
    "1111000101110001",
    "1111000110110110",
    "1111001001101101",
    "1111010000111110",
    "1111011110001100",
    "1111110000110011",
    "1111111001101000",
    "1111100101000000",
    "1111010101011000",
    "1111001101110000",
    "1111001111000010",
    "1111010111111100",
    "1111100101110010",
    "1111110101001110",
    "1111111100111101",
    "1111110011010101",
    "1111101111100100",
    "1111110010101001",
    "1111111100111010",
    "1111110001110001",
    "1111011010101000",
    "1110111111110110",
    "1110100100011010",
    "1110001011101010",
    "1101111000101100",
    "1101101101011110",
    "1101101010100101",
    "1101101111010100",
    "1101111010101010",
    "1110001011111010",
    "1110100010011001",
    "1110111101000101",
    "1111011010001100",
    "1111110110111010",
    "1111101111111100",
    "1111011101000101",
    "1111010010000000",
    "1111001110010111",
    "1111010000011001",
    "1111010101110001",
    "1111011100100001",
    "1111100011110011",
    "1111101011111010",
    "1111110101100111",
    "1111111110101011",
    "1111110001110100",
    "1111100101111011",
    "1111011101111000",
    "1111011100001100",
    "1111100010001000",
    "1111101111000100",
    "1111111111001001",
    "1111101011100010",
    "1111011000111100",
    "1111001001100000",
    "1110111110011111",
    "1110111000011010",
    "1110110111010110",
    "1110111011001111",
    "1111000011111100",
    "1111010001000111",
    "1111100001110000",
    "1111110100010011",
    "1111111001001000",
    "1111101000011100",
    "1111011011000001",
    "1111010001100111",
    "1111001100011011",
    "1111001010111010",
    "1111001100001111",
    "1111001111011010",
    "1111010011101001",
    "1111011000001110",
    "1111011100111111",
    "1111100010011001",
    "1111101001100000",
    "1111110011100110",
    "1111111110100111",
    "1111101101110010",
    "1111011100001100",
    "1111001101001111",
    "1111000100011000",
    "1111000100000110",
    "1111001101001110",
    "1111011110101110",
    "1111110110101000",
    "1111101101100010",
    "1111010000011100",
    "1110110100110110",
    "1110011101101000",
    "1110001101010111",
    "1110000101111110",
    "1110001000000001",
    "1110010010110011",
    "1110100100011100",
    "1110111010101101",
    "1111010011100010",
    "1111101101000110",
    "1111111010011011",
    "1111100101000101",
    "1111010100110110",
    "1111001011100001",
    "1111001010001001",
    "1111010000100110",
    "1111011101011011",
    "1111101110000001",
    "1111111111011111",
    "1111110000110110",
    "1111100100111100",
    "1111011101101000",
    "1111011010110000",
    "1111011011100000",
    "1111011110110011",
    "1111100011011111",
    "1111101000010111",
    "1111101100001110",
    "1111101110001101",
    "1111101101111111",
    "1111101011111001",
    "1111101001000001",
    "1111100110111000",
    "1111100110111011",
    "1111101010000111",
    "1111110000100001",
    "1111111001001110",
    "1111111101010010",
    "1111110100111100",
    "1111101111001111",
    "1111101100111111",
    "1111101110001101",
    "1111110010010000",
    "1111111000001111",
    "1111111111010111",
    "1111111000111100",
    "1111110001010010",
    "1111101010010010",
    "1111100100111001",
    "1111100010001010",
    "1111100010111001",
    "1111100111011001",
    "1111101111010110",
    "1111111001110100",
    "1111111010001110",
    "1111101101110010",
    "1111100001011110",
    "1111010101101010",
    "1111001010101111",
    "1111000001010010",
    "1110111010010011",
    "1110110111000110",
    "1110111000111111",
    "1111000001001010",
    "1111010000001010",
    "1111100101011111",
    "1111111111010101",
    "1111100101010010",
    "1111001011110111",
    "1110110111100011",
    "1110101010011011",
    "1110100101000110",
    "1110100110110010",
    "1110101110000010",
    "1110111001001110",
    "1111000111001011",
    "1111010111001000",
    "1111101000011101",
    "1111111010010111",
    "1111110100100001",
    "1111100110001000",
    "1111011100010110",
    "1111011000110100",
    "1111011100010100",
    "1111100110101000",
    "1111110110010110",
    "1111110110110011",
    "1111100011110100",
    "1111010011010010",
    "1111000111010000",
    "1111000000101100",
    "1110111111101001",
    "1111000011010111",
    "1111001010111000",
    "1111010101100111",
    "1111100011011101",
    "1111110100101000",
    "1111110111000111",
    "1111100001000101",
    "1111001011011101",
    "1110111001000110",
    "1110101100110000",
    "1110101000010101",
    "1110101100100101",
    "1110111000111010",
    "1111001011101011",
    "1111100010100111",
    "1111111011000110",
    "1111101101011101",
    "1111011001011000",
    "1111001010001111",
    "1111000000111011",
    "1110111101010111",
    "1110111110110110",
    "1111000100001011",
    "1111001100000010",
    "1111010101010111",
    "1111011111010001",
    "1111101001010011",
    "1111110011001011",
    "1111111100110100",
    "1111111001110100",
    "1111110000111001",
    "1111101000011011",
    "1111100000100011",
    "1111011001101101",
    "1111010100101001",
    "1111010010011010",
    "1111010100001010",
    "1111011010100110",
    "1111100101110111",
    "1111110101000000",
    "1111111001111001",
    "1111101001011001",
    "1111011100000001",
    "1111010011101010",
    "1111010001000101",
    "1111010011111000",
    "1111011010101010",
    "1111100011111000",
    "1111101110101000",
    "1111111010110101",
    "1111110111010110",
    "1111101000010100",
    "1111011001100000",
    "1111001101100000",
    "1111000111010000",
    "1111001000111111",
    "1111010011000011",
    "1111100011011000",
    "1111110110001100",
    "1111111000111000",
    "1111101101100000",
    "1111101001011110",
    "1111101100101100",
    "1111110101110000",
    "1111111101000110",
    "1111101101001100",
    "1111011011001001",
    "1111000111011000",
    "1110110010110001",
    "1110011110110001",
    "1110001101010010",
    "1101111111111011",
    "1101110111100011",
    "1101110011110001",
    "1101110011001111",
    "1101110100010010",
    "1101110101101001",
    "1101110110101010",
    "1101110111011111",
    "1101111000100101",
    "1101111010100110",
    "1101111101111000",
    "1110000010010111",
    "1110000111101100",
    "1110001101100000",
    "1110010011101100",
    "1110011010101000",
    "1110100011000001",
    "1110101101100001",
    "1110111010011001",
    "1111001001001100",
    "1111011000111100",
    "1111101000001110",
    "1111110101100000",
    "1111111111011010",
    "1111111010111110",
    "1111111001111111",
    "1111111101010011",
    "1111111011110011",
    "1111110010001110",
    "1111100110100010",
    "1111011001011000",
    "1111001011011101",
    "1110111101111010",
    "1110110010000110",
    "1110101001011011",
    "1110100100110111",
    "1110100100110111",
    "1110101001000010",
    "1110110000011111",
    "1110111010000111",
    "1111000100110110",
    "1111001111101100",
    "1111011001110100",
    "1111100010011010",
    "1111101000101111",
    "1111101100011000",
    "1111101101011001",
    "1111101100100010",
    "1111101011001001",
    "1111101010111101",
    "1111101101100011",
    "1111110011111011",
    "1111111110001001",
    "1111110100101111",
    "1111100110010000",
    "1111011000000001",
    "1111001011001110",
    "1111000000100100",
    "1110111000000100",
    "1110110001011010",
    "1110101100000111",
    "1110100111101101",
    "1110100100000000",
    "1110100000111101",
    "1110011110111000",
    "1110011110001100",
    "1110011111011100",
    "1110100011001011",
    "1110101001110010",
    "1110110011010111",
    "1110111111100001",
    "1111001101010110",
    "1111011011100001",
    "1111101000011111",
    "1111110011000010",
    "1111111010101011",
    "1111111111111001",
    "1111111100000010",
    "1111110111111110",
    "1111110011010000",
    "1111101110001100",
    "1111101001110010",
    "1111100111001011",
    "1111100111000011",
    "1111101001001111",
    "1111101100101111",
    "1111110000001101",
    "1111110010101010",
    "1111110011111010",
    "1111110100100010",
    "1111110101010110",
    "1111110110101101",
    "1111111000010001",
    "1111111001000101",
    "1111111000000000",
    "1111110100011001",
    "1111101110011100",
    "1111100111010010",
    "1111100000100111",
    "1111011100001001",
    "1111011011000010",
    "1111011110000000",
    "1111100101000101",
    "1111101111110110",
    "1111111101010111",
    "1111110011110111",
    "1111100101110111",
    "1111011010111010",
    "1111010101010011",
    "1111010110110010",
    "1111011111111011",
    "1111101111101111",
    "1111111100011010",
    "1111101000011000",
    "1111011000000100",
    "1111001110101000",
    "1111001101110111",
    "1111010110000110",
    "1111100110101011",
    "1111111110001001",
    "1111100101101010",
    "1111000111101000",
    "1110101010111100",
    "1110010010100001",
    "1110000000100111",
    "1101110110001001",
    "1101110010101001",
    "1101110100011101",
    "1101111001100011",
    "1110000000010010",
    "1110000111111010",
    "1110010000011110",
    "1110011010011110",
    "1110100110101000",
    "1110110101011011",
    "1111000110111011",
    "1111011010101011",
    "1111101111110111",
    "1111111010101001",
    "1111100110011010",
    "1111010101000001",
    "1111001000000001",
    "1111000000100001",
    "1110111110110000",
    "1111000001111101",
    "1111001000011000",
    "1111001111111000",
    "1111010110100010",
    "1111011011000001",
    "1111011100110111",
    "1111011100010111",
    "1111011010010100",
    "1111011000100011",
    "1111011010011001",
    "1111100011010111",
    "1111110101100010",
    "1111101111101011",
    "1111010000001010",
    "1110110001101011",
    "1110011010000111",
    "1110001101111101",
    "1110001110011110",
    "1110011001111100",
    "1110101100110010",
    "1111000010100100",
    "1111010111010011",
    "1111101000000000",
    "1111110010101111",
    "1111110110110100",
    "1111110100100110",
    "1111101100111110",
    "1111100001011010",
    "1111010011011100",
    "1111000100011111",
    "1110110110001101",
    "1110101010011110",
    "1110100011000011",
    "1110100001001101",
    "1110100101001101",
    "1110101110101001",
    "1110111100100011",
    "1111001101100110",
    "1111100000010010",
    "1111110011001111",
    "1111111010110011",
    "1111101011000010",
    "1111011110001101",
    "1111010100110001",
    "1111001110110001",
    "1111001100000001",
    "1111001100000111",
    "1111001110111000",
    "1111010100100101",
    "1111011101111111",
    "1111101011111010",
    "1111111110110100",
    "1111101001110111",
    "1111010000010010",
    "1110110111101100",
    "1110100011101010",
    "1110010111001011",
    "1110010011100100",
    "1110011000010110",
    "1110100011100001",
    "1110110010001010",
    "1111000001010010",
    "1111001110010111",
    "1111010111110010",
    "1111011100111111",
    "1111011110001111",
    "1111011100100011",
    "1111011001000100",
    "1111010100111100",
    "1111010001000111",
    "1111001110000111",
    "1111001100000111",
    "1111001010110111",
    "1111001001111100",
    "1111001000110101",
    "1111000111001011",
    "1111000100101110",
    "1111000001100100",
    "1110111110001101",
    "1110111011010001",
    "1110111001011001",
    "1110111001110100",
    "1110111110001100",
    "1111001000000110",
    "1111011000000011",
    "1111101100110100",
    "1111111100101000",
    "1111101000101101",
    "1111011011111101",
    "1111011010000110",
    "1111100100110011",
    "1111111011001000",
    "1111100110100000",
    "1111000101101100",
    "1110101000010110",
    "1110010011100100",
    "1110001010001111",
    "1110001100110011",
    "1110011001011110",
    "1110101101011100",
    "1111000110010110",
    "1111100011000011",
    "1111111100111001",
    "1111011010100101",
    "1110111000010110",
    "1110011001101010",
    "1110000010001010",
    "1101110100011000",
    "1101110001000010",
    "1101110110010011",
    "1110000000101011",
    "1110001011111100",
    "1110010100111110",
    "1110011010100101",
    "1110011101101001",
    "1110100000101001",
    "1110100110000100",
    "1110101111101001",
    "1110111101101000",
    "1111001110101001",
    "1111100000100110",
    "1111110001001100",
    "1111111110101000",
    "1111111000000101",
    "1111110011001100",
    "1111110010001111",
    "1111110100001000",
    "1111110111100001",
    "1111111011000000",
    "1111111101101101",
    "1111111111011101",
    "1111111111000110",
    "1111111101000100",
    "1111111001010001",
    "1111110011000011",
    "1111101010010111",
    "1111100000000000",
    "1111010101101110",
    "1111001101100001",
    "1111001001010101",
    "1111001010000100",
    "1111001111100011",
    "1111011000011000",
    "1111100010100100",
    "1111101011111001",
    "1111110010100101",
    "1111110101100111",
    "1111110100100101",
    "1111101111011100",
    "1111100110011000",
    "1111011001100011",
    "1111001001000110",
    "1110110101100100",
    "1110100000011110",
    "1110001100001100",
    "1101111011101000",
    "1101110001010111",
    "1101101110111111",
    "1101110100011100",
    "1110000000001000",
    "1110001111100110",
    "1110100000100100",
    "1110110010000011",
    "1111000100010010",
    "1111010111110001",
    "1111101100011001",
    "1111111111001000",
    "1111101101011010",
    "1111100001010100",
    "1111011101000100",
    "1111100001010010",
    "1111101100100111",
    "1111111100000111",
    "1111110011100001",
    "1111100101010010",
    "1111011011000001",
    "1111010101101001",
    "1111010101011010",
    "1111011010001011",
    "1111100011011100",
    "1111110000010010",
    "1111111111011010",
    "1111110000110110",
    "1111100010001010",
    "1111010101110001",
    "1111001100010110",
    "1111000101111011",
    "1111000010001111",
    "1111000001010000",
    "1111000011011100",
    "1111001001011101",
    "1111010011111100",
    "1111100011000011",
    "1111110101110010",
    "1111110101110000",
    "1111100010011100",
    "1111010011001011",
    "1111001010010011",
    "1111001001001011",
    "1111001111110001",
    "1111011100111111",
    "1111101110101000",
    "1111111101110010",
    "1111101010111100",
    "1111011010111010",
    "1111001111000111",
    "1111001000001011",
    "1111000110000011",
    "1111001000001000",
    "1111001101100000",
    "1111010101001110",
    "1111011110101101",
    "1111101001111011",
    "1111110111110111",
    "1111110101111000",
    "1111011110010110",
    "1111000010001000",
    "1110100100000001",
    "1110001000100010",
    "1101110100011111",
    "1101101011011001",
    "1101101110001111",
    "1101111010111101",
    "1110001101010111",
    "1110100000110000",
    "1110110001101011",
    "1110111111111011",
    "1111001110101110",
    "1111100010001010",
    "1111111100010111",
    "1111100100000110",
    "1111000100100101",
    "1110101011111100",
    "1110100000001101",
    "1110100100011000",
    "1110110110101111",
    "1111010010010101",
    "1111110001001000",
    "1111110010001111",
    "1111011011010110",
    "1111001100000010",
    "1111000101000110",
    "1111000110011101",
    "1111001111100001",
    "1111011111010111",
    "1111110100001011",
    "1111110100101011",
    "1111011110011100",
    "1111001100011011",
    "1111000001000000",
    "1110111101001100",
    "1111000000001101",
    "1111000111111111",
    "1111010010010010",
    "1111011101001100",
    "1111100111010010",
    "1111101111101101",
    "1111110101111101",
    "1111111001111111",
    "1111111100010000",
    "1111111101110000",
    "1111111111110000",
    "1111111100011101",
    "1111110110000110",
    "1111101101000110",
    "1111100010010100",
    "1111010111010101",
    "1111001110001010",
    "1111001000100101",
    "1111000111110101",
    "1111001100010100",
    "1111010101011010",
    "1111100010001010",
    "1111110001100101",
    "1111111101010001",
    "1111101011100110",
    "1111011011000110",
    "1111001101110000",
    "1111000101010111",
    "1111000010101110",
    "1111000101011011",
    "1111001100000100",
    "1111010100110110",
    "1111011110010001",
    "1111100111111100",
    "1111110010011110",
    "1111111111001010",
    "1111110000111100",
    "1111011110000101",
    "1111001010000110",
    "1110111000001000",
    "1110101011101111",
    "1110100111110100",
    "1110101101101011",
    "1110111100110011",
    "1111010011001000",
    "1111101101011010",
    "1111110111111000",
    "1111100000001100",
    "1111001110010100",
    "1111000100010010",
    "1111000011001000",
    "1111001010101011",
    "1111011001100011",
    "1111101101001110",
    "1111111101100100",
    "1111101010011000",
    "1111011100001110",
    "1111010101010000",
    "1111010110010000",
    "1111011110101110",
    "1111101101011011",
    "1111111111010101",
    "1111101001101101",
    "1111010011111110",
    "1111000000100001",
    "1110110001010000",
    "1110100111011000",
    "1110100010110011",
    "1110100010011100",
    "1110100100110011",
    "1110101000101111",
    "1110101110010110",
    "1110110110110001",
    "1111000011101100",
    "1111010110011010",
    "1111101110110001",
    "1111110101001101",
    "1111011000111111",
    "1111000000100111",
    "1110101111011001",
    "1110100110111100",
    "1110100111000001",
    "1110101101111010",
    "1110111001010001",
    "1111000110111110",
    "1111010101100101",
    "1111100100001101",
    "1111110010001010",
    "1111111110100111",
    "1111110111011000",
    "1111110000101110",
    "1111101101110101",
    "1111101110101000",
    "1111110010101000",
    "1111111001000011",
    "1111111110101001",
    "1111110100111010",
    "1111101001111000",
    "1111011101110011",
    "1111010001011001",
    "1111000101101111",
    "1110111100001111",
    "1110110110000100",
    "1110110011111001",
    "1110110101101001",
    "1110111010110101",
    "1111000011000110",
    "1111001110100100",
    "1111011101111000",
    "1111110001100001",
    "1111110110111110",
    "1111011101110010",
    "1111000110011101",
    "1110110101001000",
    "1110101101001100",
    "1110110000001000",
    "1110111101000101",
    "1111010001001101",
    "1111101000100101",
    "1111111111010000",
    "1111101110000110",
    "1111100010000101",
    "1111011110011011",
    "1111100100000011",
    "1111110010111101",
    "1111110110010000",
    "1111011010011101",
    "1110111101011001",
    "1110100011000000",
    "1110001110011011",
    "1110000001010101",
    "1101111011110101",
    "1101111100101010",
    "1110000010010100",
    "1110001011110000",
    "1110011000101101",
    "1110101001001011",
    "1110111100110000",
    "1111010010010101",
    "1111100111110010",
    "1111111010100100",
    "1111110111010000",
    "1111101110100110",
    "1111101010100110",
    "1111101001010111",
    "1111101000100111",
    "1111100110100000",
    "1111100010010000",
    "1111011100010011",
    "1111010101101111",
    "1111010000000010",
    "1111001100010110",
    "1111001011000010",
    "1111001011110101",
    "1111001101110111",
    "1111010000000011",
    "1111010001100110",
    "1111010010001111",
    "1111010010101110",
    "1111010101000001",
    "1111011011101101",
    "1111101000100011",
    "1111111011101000",
    "1111101101000100",
    "1111010101011101",
    "1111000010000010",
    "1110110110011011",
    "1110110100010010",
    "1110111010101101",
    "1111000111000011",
    "1111010101111011",
    "1111100100001010",
    "1111101111101010",
    "1111110111000111",
    "1111111001111001",
    "1111110111101111",
    "1111110000101101",
    "1111100101010010",
    "1111010110101111",
    "1111000111000001",
    "1110111000100010",
    "1110101101110000",
    "1110101000011110",
    "1110101001101011",
    "1110110001011110",
    "1110111111011001",
    "1111010010100001",
    "1111101001010000",
    "1111111110101100",
    "1111101000011010",
    "1111010110101100",
    "1111001011100000",
    "1111000111010101",
    "1111001000111100",
    "1111001110000100",
    "1111010100000001",
    "1111011000111001",
    "1111011100000010",
    "1111011110010100",
    "1111100001100111",
    "1111101000001000",
    "1111110011010010",
    "1111111100111001",
    "1111101010000011",
    "1111010111000001",
    "1111000111001000",
    "1110111101001001",
    "1110111010101010",
    "1110111111110000",
    "1111001011001110",
    "1111011010110111",
    "1111101100000100",
    "1111111100010100",
    "1111110110011010",
    "1111101101010101",
    "1111101000100111",
    "1111100111101111",
    "1111101001101011",
    "1111101101010111",
    "1111110001110110",
    "1111110110101011",
    "1111111011110011",
    "1111111110011001",
    "1111110111100001",
    "1111101110111101",
    "1111100100011101",
    "1111011000010011",
    "1111001011100011",
    "1110111111110110",
    "1110110111000001",
    "1110110010100010",
    "1110110011011010",
    "1110111001101111",
    "1111000101000101",
    "1111010100011101",
    "1111100110101011",
    "1111111010000010",
    "1111110011011010",
    "1111100011111011",
    "1111011001100011",
    "1111010101110100",
    "1111011001010000",
    "1111100011000101",
    "1111110001011011",
    "1111111110010111",
    "1111101111001000",
    "1111100011010101",
    "1111011100111000",
    "1111011100111111",
    "1111100011111100",
    "1111110001001111",
    "1111111100101100",
    "1111101000010110",
    "1111010100101100",
    "1111000100110011",
    "1110111011010100",
    "1110111001111111",
    "1111000001100100",
    "1111010001011111",
    "1111100111110101",
    "1111111110011000",
    "1111100100110100",
    "1111001110101000",
    "1110111101111111",
    "1110110011100100",
    "1110101110100100",
    "1110101101001010",
    "1110101101001111",
    "1110101101000111",
    "1110101100000010",
    "1110101010000100",
    "1110100111101111",
    "1110100101110111",
    "1110100101000101",
    "1110100101110010",
    "1110101000000011",
    "1110101011101010",
    "1110110000010010",
    "1110110101011101",
    "1110111010111000",
    "1111000001001111",
    "1111001010010100",
    "1111011000010011",
    "1111101100011111",
    "1111111001101101",
    "1111011101001010",
    "1111000010000000",
    "1110101100011011",
    "1110011111001111",
    "1110011010101011",
    "1110011101001010",
    "1110100100011101",
    "1110101111001100",
    "1110111101001001",
    "1111001110101000",
    "1111100011001010",
    "1111111000110011",
    "1111110011100101",
    "1111100101101010",
    "1111100000000000",
    "1111100011001111",
    "1111101110000101",
    "1111111110001101",
    "1111101111000100",
    "1111011100000001",
    "1111001010001110",
    "1110111010111100",
    "1110101111010110",
    "1110101000110101",
    "1110101000110100",
    "1110110000010111",
    "1110111111110011",
    "1111010110000110",
    "1111110000101111",
    "1111110100001010",
    "1111011100111100",
    "1111001101000111",
    "1111000110011111",
    "1111001000101010",
    "1111010001010101",
    "1111011101010001",
    "1111101001001101",
    "1111110011000000",
    "1111111001111111",
    "1111111110100100",
    "1111111110010000",
    "1111111011101000",
    "1111111001000100",
    "1111110110101011",
    "1111110101001001",
    "1111110101011011",
    "1111111000010011",
    "1111111110001101",
    "1111111001000001",
    "1111101110000100",
    "1111100010000011",
    "1111010110011010",
    "1111001100101000",
    "1111000110000100",
    "1111000011100100",
    "1111000101011000",
    "1111001011011001",
    "1111010101010000",
    "1111100010100001",
    "1111110010100111",
    "1111111011010001",
    "1111101000011011",
    "1111010110000011",
    "1111000101000110",
    "1110110110000110",
    "1110101001001011",
    "1110011110001101",
    "1110010101000011",
    "1110001101100110",
    "1110000111101101",
    "1110000011001011",
    "1101111111110000",
    "1101111101000010",
    "1101111010110111",
    "1101111001001011",
    "1101110111111110",
    "1101110111010000",
    "1101110110110010",
    "1101110110001001",
    "1101110100111110",
    "1101110011001000",
    "1101110001000000",
    "1101101111011001",
    "1101101111010001",
    "1101110001011111",
    "1101110110011101",
    "1101111101111010",
    "1110000111000001",
    "1110010000110011",
    "1110011010011000",
    "1110100011010010",
    "1110101100100101",
    "1110111001010000",
    "1111001100010011",
    "1111100110101000",
    "1111111010000011",
    "1111011011001110",
    "1111000010111110",
    "1110110110010110",
    "1110110111011111",
    "1111000100010101",
    "1111011000000011",
    "1111101101010010",
    "1111111111110110",
    "1111110000110111",
    "1111100101001011",
    "1111011011110101",
    "1111010100000001",
    "1111001101111000",
    "1111001010011011",
    "1111001010101010",
    "1111001110111111",
    "1111010110110111",
    "1111100000111011",
    "1111101011011010",
    "1111110101001110",
    "1111111110001111",
    "1111111000111010",
    "1111101111110010",
    "1111100110001110",
    "1111011100101101",
    "1111010011101110",
    "1111001100000001",
    "1111000110001101",
    "1111000010111001",
    "1111000010110100",
    "1111000110110110",
    "1111001111111000",
    "1111011110110101",
    "1111110011101111",
    "1111110010101100",
    "1111010111100010",
    "1110111110110001",
    "1110101100010100",
    "1110100010101111",
    "1110100010100001",
    "1110101001110010",
    "1110110101100111",
    "1111000011100010",
    "1111010010110100",
    "1111100100011000",
    "1111111001001001",
    "1111101111001101",
    "1111010111001011",
    "1111000010011111",
    "1110110100101100",
    "1110101111110101",
    "1110110011101100",
    "1110111110001100",
    "1111001100101110",
    "1111011101101001",
    "1111110000101110",
    "1111111001110101",
    "1111100010111101",
    "1111001101000101",
    "1110111100001010",
    "1110110100000011",
    "1110110110111011",
    "1111000100010010",
    "1111011001010110",
    "1111110010010001",
    "1111110100000001",
    "1111011011000100",
    "1111000011001010",
    "1110101100100001",
    "1110011000010101",
    "1110001001000110",
    "1110000010001010",
    "1110000110010101",
    "1110010110100000",
    "1110110000111000",
    "1111010001010010",
    "1111110010010010",
    "1111110001001001",
    "1111011100010110",
    "1111010000000101",
    "1111001011001100",
    "1111001011010110",
    "1111001110010001",
    "1111010010011100",
    "1111010111001101",
    "1111011100110000",
    "1111100011100010",
    "1111101011110001",
    "1111110101010000",
    "1111111111011000",
    "1111110110110000",
    "1111101110010100",
    "1111101000011001",
    "1111100101111011",
    "1111100111011010",
    "1111101100101010",
    "1111110100101101",
    "1111111101111100",
    "1111111001011110",
    "1111110011010111",
    "1111110000111100",
    "1111110010100101",
    "1111110111111110",
    "1111111111101001",
    "1111110101000110",
    "1111101000111001",
    "1111011011100000",
    "1111001101011011",
    "1110111111011100",
    "1110110010101001",
    "1110101000000100",
    "1110100000101100",
    "1110011101001001",
    "1110011101101000",
    "1110100010000110",
    "1110101010101010",
    "1110110111011111",
    "1111001000111110",
    "1111011110111111",
    "1111111000010110",
    "1111101101100000",
    "1111010110001101",
    "1111000101001110",
    "1110111101001010",
    "1110111110011111",
    "1111000111101000",
    "1111010101011000",
    "1111100100011010",
    "1111110010111110",
    "1111111110001001",
    "1111101100101111",
    "1111010110101100",
    "1110111100000010",
    "1110011111100100",
    "1110000110001001",
    "1101110101000011",
    "1101101111111111",
    "1101110111101000",
    "1110001001101111",
    "1110100010001111",
    "1110111100101101",
    "1111010101011011",
    "1111101001110011",
    "1111111000001010",
    "1111111111100100",
    "1111111111101100",
    "1111111000101111",
    "1111101011101110",
    "1111011010100011",
    "1111000111111100",
    "1110110111001000",
    "1110101010111111",
    "1110100101100100",
    "1110100111011101",
    "1110110000000000",
    "1110111101100011",
    "1111001110000000",
    "1111011111010001",
    "1111101111011001",
    "1111111101000011",
    "1111111000011110",
    "1111110001000111",
    "1111101011111000",
    "1111100111010111",
    "1111100010001010",
    "1111011011011011",
    "1111010011010010",
    "1111001010101011",
    "1111000011010010",
    "1110111110110000",
    "1110111110001111",
    "1111000010000110",
    "1111001001110000",
    "1111010100000101",
    "1111011111111011",
    "1111101101000001",
    "1111111011111010",
    "1111110010011110",
    "1111011110000010",
    "1111001000001011",
    "1110110011111011",
    "1110100100101111",
    "1110011101010110",
    "1110011110011100",
    "1110100110100101",
    "1110110010101110",
    "1110111111010001",
    "1111001001010101",
    "1111001111101100",
    "1111010010101001",
    "1111010011010101",
    "1111010011001010",
    "1111010011000011",
    "1111010011011000",
    "1111010100000000",
    "1111010100001101",
    "1111010011010010",
    "1111010000100100",
    "1111001011101111",
    "1111000100111001",
    "1110111100101010",
    "1110110100010010",
    "1110101101100011",
    "1110101010100101",
    "1110101101000100",
    "1110110101110010",
    "1111000100001101",
    "1111010110100000",
    "1111101001111100",
    "1111111011010100",
    "1111111000001000",
    "1111110010011001",
    "1111110011111101",
    "1111111100001001",
    "1111110110101111",
    "1111100111000010",
    "1111010111001101",
    "1111001001100010",
    "1110111111110000",
    "1110111010111100",
    "1110111011001110",
    "1111000000001000",
    "1111001000101100",
    "1111010011110001",
    "1111100000101001",
    "1111101111000100",
    "1111111111001001",
    "1111101111000011",
    "1111011100000010",
    "1111001000111001",
    "1110110110111110",
    "1110100111101000",
    "1110011011101010",
    "1110010011001000",
    "1110001101011110",
    "1110001010000010",
    "1110001000100011",
    "1110001001011001",
    "1110001101100100",
    "1110010110001001",
    "1110100011111000",
    "1110110110011111",
    "1111001100110011",
    "1111100100110110",
    "1111111011111101",
    "1111110000011111",
    "1111100010101110",
    "1111011011110010",
    "1111011011100000",
    "1111100000011100",
    "1111101000100001",
    "1111110001100000",
    "1111111001111100",
    "1111111110011111",
    "1111110110111001",
    "1111101101100101",
    "1111100001010010",
    "1111010001111110",
    "1111000001010100",
    "1110110001111011",
    "1110100110101101",
    "1110100001100010",
    "1110100010111101",
    "1110101001111111",
    "1110110100110001",
    "1111000001010000",
    "1111001101101000",
    "1111011000010001",
    "1111011111101001",
    "1111100010001000",
    "1111011110010111",
    "1111010011110110",
    "1111000011011101",
    "1110101111011100",
    "1110011011001100",
    "1110001010011011",
    "1110000000001100",
    "1101111110010110",
    "1110000101010000",
    "1110010100000011",
    "1110101001000010",
    "1111000010001000",
    "1111011100111010",
    "1111110110111111",
    "1111110001111001",
    "1111011111101011",
    "1111010011010111",
    "1111001100110101",
    "1111001010111100",
    "1111001011101010",
    "1111001100111101",
    "1111001101010001",
    "1111001011110101",
    "1111001000111110",
    "1111000101100100",
    "1111000010110110",
    "1111000001111000",
    "1111000011010111",
    "1111000111100111",
    "1111001110011111",
    "1111010111110001",
    "1111100011001000",
    "1111110000011001",
    "1111111111010001",
    "1111110000100011",
    "1111011111111010",
    "1111001111111101",
    "1111000010001011",
    "1110110111111110",
    "1110110010000000",
    "1110110000010010",
    "1110110010000101",
    "1110110110010110",
    "1110111100010110",
    "1111000100000011",
    "1111001110000111",
    "1111011011010100",
    "1111101011111010",
    "1111111110111001",
    "1111101101110100",
    "1111011101000100",
    "1111010001010111",
    "1111001100000001",
    "1111001100111010",
    "1111010010100001",
    "1111011010101010",
    "1111100011000011",
    "1111101010000110",
    "1111101110111010",
    "1111110001001000",
    "1111110000101100",
    "1111101101101011",
    "1111101000011000",
    "1111100001100010",
    "1111011010010110",
    "1111010100010000",
    "1111010000101110",
    "1111010000101100",
    "1111010100011101",
    "1111011011100000",
    "1111100100110011",
    "1111101111000011",
    "1111111001001010",
    "1111111101100110",
    "1111110101101100",
    "1111101111010110",
    "1111101010101110",
    "1111100111111110",
    "1111100111001010",
    "1111101000001110",
    "1111101010111110",
    "1111101111001010",
    "1111110100100011",
    "1111111011001001",
    "1111111101000110",
    "1111110100010101",
    "1111101010111001",
    "1111100001100001",
    "1111011001001100",
    "1111010011000011",
    "1111010000000010",
    "1111010000101100",
    "1111010101001101",
    "1111011101001111",
    "1111101000000110",
    "1111110100111101",
    "1111111100111100",
    "1111101110001111",
    "1111011111010110",
    "1111010000100011",
    "1111000010010100",
    "1110110101010000",
    "1110101010000111",
    "1110100001100111",
    "1110011100000111",
    "1110011001100010",
    "1110011001011000",
    "1110011010111111",
    "1110011101111010",
    "1110100010000011",
    "1110100111101101",
    "1110101111010010",
    "1110111000101000",
    "1111000010111011",
    "1111001100101101",
    "1111010100000110",
    "1111010111101101",
    "1111010110111001",
    "1111010010010101",
    "1111001011110010",
    "1111000101101010",
    "1111000010011111",
    "1111000100010010",
    "1111001100011100",
    "1111011011011101",
    "1111110000101111",
    "1111110101011101",
    "1111011010000111",
    "1111000000101110",
    "1110101100100000",
    "1110011111101100",
    "1110011011000111",
    "1110011101111111",
    "1110100110100000",
    "1110110010101001",
    "1111000000111110",
    "1111010000111110",
    "1111100010100110",
    "1111110101100010",
    "1111110111001010",
    "1111100101100000",
    "1111010111111001",
    "1111010000011111",
    "1111010000010111",
    "1111010110111110",
    "1111100010010000",
    "1111101111010100",
    "1111111011010110",
    "1111111011100110",
    "1111110110011101",
    "1111110101000100",
    "1111110110101000",
    "1111111010000011",
    "1111111110001100",
    "1111111101111101",
    "1111111011011101",
    "1111111011000001",
    "1111111101001101",
    "1111111101111010",
    "1111110111000011",
    "1111101111011010",
    "1111101000101110",
    "1111100100101010",
    "1111100100101110",
    "1111101001100111",
    "1111110011010011",
    "1111111111001000",
    "1111101111100011",
    "1111011111111010",
    "1111010010000011",
    "1111000111010001",
    "1111000000000111",
    "1110111100011011",
    "1110111011101010",
    "1110111101010100",
    "1111000001011001",
    "1111001000011010",
    "1111010011001010",
    "1111100010000110",
    "1111110100100010",
    "1111110111011111",
    "1111100100111011",
    "1111010110110001",
    "1111001111000111",
    "1111001110101000",
    "1111010100101001",
    "1111011111101001",
    "1111101110000111",
    "1111111110100111",
    "1111110000010011",
    "1111100000011111",
    "1111010011110001",
    "1111001011110111",
    "1111001001111100",
    "1111001110011001",
    "1111011000110100",
    "1111101000011000",
    "1111111100000100",
    "1111101101010001",
    "1111010101011010",
    "1110111110101000",
    "1110101011100011",
    "1110011110100110",
    "1110011001011000",
    "1110011100001110",
    "1110100110001101",
    "1110110101100100",
    "1111001000011110",
    "1111011101101000",
    "1111110100010000",
    "1111110100010100",
    "1111011101001100",
    "1111000111111111",
    "1110110110101100",
    "1110101011000001",
    "1110100101110100",
    "1110100110110001",
    "1110101100010111",
    "1110110100111011",
    "1110111111000010",
    "1111001010001011",
    "1111010110100101",
    "1111100100110001",
    "1111110100111010",
    "1111111001101011",
    "1111101000100101",
    "1111011001110101",
    "1111001111010010",
    "1111001010000100",
    "1111001010010001",
    "1111001111000000",
    "1111010110110001",
    "1111100000000010",
    "1111101001101001",
    "1111110010111101",
    "1111111011011100",
    "1111111101011111",
    "1111111000101101",
    "1111110110111111",
    "1111111000111101",
    "1111111110110000",
    "1111110111111110",
    "1111101100000111",
    "1111011110110101",
    "1111010001100001",
    "1111000101110010",
    "1110111101010110",
    "1110111001111101",
    "1110111101000111",
    "1111000111101100",
    "1111011001001100",
    "1111101111101110",
    "1111110111111111",
    "1111100001110011",
    "1111010000111011",
    "1111000111011010",
    "1111000101011111",
    "1111001001110100",
    "1111010010000000",
    "1111011011110111",
    "1111100110011000",
    "1111110010001000",
    "1111111111011101",
    "1111101101011001",
    "1111011000000011",
    "1111000001100100",
    "1110101101100100",
    "1110100000000010",
    "1110011011111010",
    "1110100001111110",
    "1110110000101100",
    "1111000100101001",
    "1111011001100011",
    "1111101011100011",
    "1111110111101111",
    "1111111100100100",
    "1111111001110110",
    "1111110000100111",
    "1111100010110011",
    "1111010010111001",
    "1111000011011101",
    "1110110110101100",
    "1110101110000000",
    "1110101001111100",
    "1110101010000010",
    "1110101101001111",
    "1110110010001101",
    "1110110111110010",
    "1110111101001111",
    "1111000010000010",
    "1111000101111011",
    "1111001000110100",
    "1111001010111000",
    "1111001100100000",
    "1111001110011100",
    "1111010001110110",
    "1111010111111110",
    "1111100001111000",
    "1111101111101110",
    "1111111111100000",
    "1111101110001011",
    "1111011111000000",
    "1111010100011111",
    "1111001111111011",
    "1111010001010000",
    "1111010111000110",
    "1111011111011111",
    "1111101000111111",
    "1111110011001101",
    "1111111110111001",
    "1111110011000000",
    "1111100010011111",
    "1111010000111011",
    "1111000001000000",
    "1110110101101010",
    "1110110001000000",
    "1110110011010010",
    "1110111011000110",
    "1111000110001001",
    "1111010010011101",
    "1111011111011111",
    "1111101101111111",
    "1111111110111111",
    "1111101101011110",
    "1111011001010001",
    "1111000111100101",
    "1110111011111111",
    "1110111001000111",
    "1110111111110110",
    "1111001111001000",
    "1111100100011101",
    "1111111100111110",
    "1111101001111010",
    "1111010010011101",
    "1110111110101001",
    "1110110000010111",
    "1110101001100000",
    "1110101011100001",
    "1110110110111011",
    "1111001010100110",
    "1111100011111000",
    "1111111111000000",
    "1111100111110010",
    "1111010011011101",
    "1111000101010011",
    "1110111101001010",
    "1110111001110101",
    "1110111001111111",
    "1110111100111010",
    "1111000010101001",
    "1111001011111000",
    "1111011001010110",
    "1111101011000111",
    "1111111111101100",
    "1111101001001011",
    "1111010100000001",
    "1111000011000101",
    "1110111000100011",
    "1110110101100101",
    "1110111010001001",
    "1111000100111110",
    "1111010100000110",
    "1111100101000101",
    "1111110101100001",
    "1111111100101101",
    "1111110011001110",
    "1111101110110111",
    "1111101111101011",
    "1111110101000100",
    "1111111110000100",
    "1111110110010111",
    "1111101001010110",
    "1111011011110101",
    "1111001110110101",
    "1111000011010011",
    "1110111010001110",
    "1110110100010000",
    "1110110001110001",
    "1110110010101111",
    "1110110110101010",
    "1110111100110010",
    "1111000100100101",
    "1111001110111000",
    "1111011101100100",
    "1111110010100011",
    "1111110001111010",
    "1111010010001011",
    "1110110010110001",
    "1110011000111100",
    "1110001001001011",
    "1110000101010011",
    "1110001011110111",
    "1110011001000001",
    "1110101000010000",
    "1110110110110110",
    "1111000100110011",
    "1111010011111000",
    "1111100101101110",
    "1111111010010101",
    "1111110000101111",
    "1111011111110110",
    "1111010111101010",
    "1111011011001110",
    "1111101010011001",
    "1111111110010000",
    "1111100100011000",
    "1111001101110000",
    "1110111110110001",
    "1110111001110010",
    "1110111111010010",
    "1111001101111111",
    "1111100011001111",
    "1111111011011101",
    "1111101101000111",
    "1111011001111001",
    "1111001100110111",
    "1111000110101100",
    "1111000110100010",
    "1111001010011110",
    "1111010000000111",
    "1111010101101001",
    "1111011010001100",
    "1111011101111101",
    "1111100001100100",
    "1111100101100000",
    "1111101001111010",
    "1111101110011001",
    "1111110010011011",
    "1111110101100101",
    "1111110111110100",
    "1111111001011100",
    "1111111010111001",
    "1111111100010111",
    "1111111110001001",
    "1111111110010110",
    "1111110111000111",
    "1111101010010000",
    "1111010111011010",
    "1111000000011111",
    "1110101001010000",
    "1110010110000100",
    "1110001010101101",
    "1110001000101111",
    "1110001111001101",
    "1110011011011001",
    "1110101010000100",
    "1110111000101101",
    "1111000110000100",
    "1111010001101100",
    "1111011011011000",
    "1111100010101100",
    "1111100110011110",
    "1111100101010111",
    "1111011110001001",
    "1111010000011110",
    "1110111101010110",
    "1110100111001011",
    "1110010001001010",
    "1101111110010010",
    "1101110000110001",
    "1101101001111010",
    "1101101001111001",
    "1101110000000011",
    "1101111010111000",
    "1110001000100000",
    "1110010111001101",
    "1110100101101010",
    "1110110011001000",
    "1110111111000100",
    "1111001001000001",
    "1111010000101001",
    "1111010101100100",
    "1111010111100000",
    "1111010110101000",
    "1111010011100111",
    "1111001111100110",
    "1111001100000001",
    "1111001010001111",
    "1111001011100011",
    "1111010000110000",
    "1111011010001001",
    "1111100111001111",
    "1111110110111111",
    "1111111000000110",
    "1111100111101011",
    "1111011001001001",
    "1111001101011011",
    "1111000101000011",
    "1111000000010001",
    "1110111111001000",
    "1111000001111000",
    "1111001001000010",
    "1111010101010000",
    "1111100110101111",
    "1111111100101101",
    "1111101010110010",
    "1111010010100111",
    "1110111101101011",
    "1110101110010001",
    "1110100101100000",
    "1110100011010000",
    "1110100110011011",
    "1110101101101011",
    "1110110111111111",
    "1111000100111011",
    "1111010100010000",
    "1111100101101100",
    "1111111000011110",
    "1111110100100111",
    "1111100011010010",
    "1111010101000101",
    "1111001011000111",
    "1111000101110001",
    "1111000100100111",
    "1111000110111001",
    "1111001011110101",
    "1111010010110001",
    "1111011011001100",
    "1111100100100101",
    "1111101110010010",
    "1111110111011010",
    "1111111110111011",
    "1111111100011011",
    "1111111100000001",
    "1111111111000010",
    "1111110100010000",
    "1111100100000000",
    "1111001111101110",
    "1110111001110000",
    "1110100100111011",
    "1110010011111001",
    "1110001000110010",
    "1110000100100101",
    "1110000111011111",
    "1110010000111101",
    "1110100000010010",
    "1110110100101100",
    "1111001100111010",
    "1111100111000110",
    "1111111111010101",
    "1111101001101001",
    "1111011010111100",
    "1111010101011000",
    "1111011001101010",
    "1111100110101001",
    "1111111001101111",
    "1111110000011101",
    "1111011011100011",
    "1111001010011011",
    "1110111111001000",
    "1110111010100011",
    "1110111100100011",
    "1111000011111110",
    "1111001111000100",
    "1111011011101111",
    "1111101000000100",
    "1111110010100001",
    "1111111010001101",
    "1111111110111011",
    "1111111110110010",
    "1111111110000001",
    "1111111101010110",
    "1111111011010101",
    "1111110110101111",
    "1111101110110101",
    "1111100011101100",
    "1111010110000110",
    "1111000111011111",
    "1110111001101011",
    "1110101110011110",
    "1110100111001001",
    "1110100100001101",
    "1110100101010011",
    "1110101001011011",
    "1110101111000100",
    "1110110100111001",
    "1110111010001111",
    "1110111111110000",
    "1111000111001110",
    "1111010011000001",
    "1111100100110110",
    "1111111100100011",
    "1111101000000000",
    "1111001100111101",
    "1110110110110001",
    "1110101000111111",
    "1110100101000001",
    "1110101001110010",
    "1110110100100101",
    "1111000010010111",
    "1111010000100110",
    "1111011101111101",
    "1111101010001000",
    "1111110100111111",
    "1111111110000111",
    "1111111011101001",
    "1111111001110001",
    "1111111101001000",
    "1111111010011110",
    "1111101110111011",
    "1111100011000110",
    "1111011010010011",
    "1111010111000011",
    "1111011010100101",
    "1111100100100100",
    "1111110011001001",
    "1111111100010001",
    "1111101100101010",
    "1111100000010100",
    "1111011000100000",
    "1111010101011000",
    "1111010110000110",
    "1111011001001011",
    "1111011101001110",
    "1111100001001000",
    "1111100100101010",
    "1111101000001110",
    "1111101100101111",
    "1111110011010011",
    "1111111100101101",
    "1111110110110000",
    "1111100111101011",
    "1111010111010000",
    "1111000111000110",
    "1110111000110100",
    "1110101101101110",
    "1110100110110110",
    "1110100100100100",
    "1110100110101101",
    "1110101100101010",
    "1110110101001000",
    "1110111110101011",
    "1111000111111010",
    "1111001111110110",
    "1111010110001101",
    "1111011011010110",
    "1111100000010010",
    "1111100110000110",
    "1111101101101000",
    "1111110110111111",
    "1111111110010111",
    "1111110011101110",
    "1111101010011001",
    "1111100011100111",
    "1111100000001100",
    "1111100000010100",
    "1111100011110100",
    "1111101010001111",
    "1111110010110101",
    "1111111100100010",
    "1111111001111000",
    "1111110001111101",
    "1111101100111101",
    "1111101011101110",
    "1111101110010000",
    "1111110011101100",
    "1111111010011011",
    "1111111111011011",
    "1111111011110110",
    "1111111100001010",
    "1111111110111100",
    "1111110101101010",
    "1111101000101100",
    "1111011001010001",
    "1111001001000111",
    "1110111010010001",
    "1110101110110011",
    "1110101000011110",
    "1110101000001100",
    "1110101101110010",
    "1110110111110111",
    "1111000100010000",
    "1111010000011111",
    "1111011010011101",
    "1111100000110001",
    "1111100011000101",
    "1111100001101110",
    "1111011101100100",
    "1111010111110001",
    "1111010001100010",
    "1111001100000001",
    "1111001000001001",
    "1111000110100111",
    "1111000111101111",
    "1111001011010001",
    "1111010000010010",
    "1111010101001101",
    "1111011000001000",
    "1111010111010000",
    "1111010001011111",
    "1111000110101111",
    "1110111000000100",
    "1110100111011101",
    "1110010111010011",
    "1110001001111001",
    "1110000000111101",
    "1101111101010001",
    "1101111110101011",
    "1110000100010111",
    "1110001101011100",
    "1110011001100111",
    "1110101001001100",
    "1110111100110000",
    "1111010100010111",
    "1111101111000011",
    "1111110101011111",
    "1111011100010110",
    "1111001000010101",
    "1110111011000100",
    "1110110100100010",
    "1110110011011000",
    "1110110101101010",
    "1110111001101010",
    "1110111110100011",
    "1111000100001000",
    "1111001010100101",
    "1111010001100111",
    "1111011000001011",
    "1111011100100000",
    "1111011100100011",
    "1111010110110001",
    "1111001010110111",
    "1110111010000111",
    "1110100111000110",
    "1110010100111011",
    "1110000110100100",
    "1101111110000010",
    "1101111100010011",
    "1110000001010100",
    "1110001100100011",
    "1110011101011100",
    "1110110011011101",
    "1111001101110000",
    "1111101010110110",
    "1111110111110101",
    "1111011101100100",
    "1111001001011101",
    "1110111101100001",
    "1110111010001011",
    "1110111101111111",
    "1111000110100010",
    "1111010001001111",
    "1111011100010100",
    "1111100111001100",
    "1111110010001110",
    "1111111110001001",
    "1111110100100011",
    "1111100110001101",
    "1111010111101101",
    "1111001010101010",
    "1111000000110001",
    "1110111011100011",
    "1110111011110101",
    "1111000001100111",
    "1111001100001001",
    "1111011001111010",
    "1111101000111010",
    "1111110110111100",
    "1111111101111110",
    "1111110111011101",
    "1111110110001000",
    "1111111001110010",
    "1111111110011111",
    "1111110100001010",
    "1111101000110010",
    "1111011101110101",
    "1111010100011100",
    "1111001101010010",
    "1111001000111010",
    "1111000111011011",
    "1111001000111010",
    "1111001101001110",
    "1111010100000101",
    "1111011100111111",
    "1111100111011000",
    "1111110010100100",
    "1111111101111001",
    "1111110111010100",
    "1111101101110101",
    "1111100110010010",
    "1111100001010101",
    "1111011111011111",
    "1111100001000111",
    "1111100110010010",
    "1111101111000010",
    "1111111011101011",
    "1111110011010011",
    "1111011110000010",
    "1111000101101001",
    "1110101100101011",
    "1110010110100010",
    "1110000110100101",
    "1101111111001010",
    "1110000000110110",
    "1110001010001111",
    "1110011000100111",
    "1110101001100011",
    "1110111100011100",
    "1111010010000010",
    "1111101011000111",
    "1111111000110110",
    "1111011100100011",
    "1111000100001000",
    "1110110011111011",
    "1110101110101011",
    "1110110100000000",
    "1111000000100001",
    "1111001111010111",
    "1111011011111101",
    "1111100011101010",
    "1111100110001101",
    "1111100100111001",
    "1111100001110011",
    "1111011110100110",
    "1111011100001001",
    "1111011010100010",
    "1111011001100000",
    "1111011000110111",
    "1111011000100101",
    "1111011000111001",
    "1111011001110000",
    "1111011010110101",
    "1111011011011101",
    "1111011011001111",
    "1111011010010110",
    "1111011001011011",
    "1111011001011000",
    "1111011011000010",
    "1111011111000100",
    "1111100101110110",
    "1111101111101011",
    "1111111100111010",
    "1111110010001110",
    "1111011110000000",
    "1111000111110010",
    "1110110001111011",
    "1110011111010111",
    "1110010010110100",
    "1110001101111000",
    "1110010000011001",
    "1110011000100010",
    "1110100011010011",
    "1110101101101011",
    "1110110101100010",
    "1110111010100010",
    "1110111110010001",
    "1111000011011111",
    "1111001100100110",
    "1111011010011000",
    "1111101011010011",
    "1111111100010001",
    "1111110110011110",
    "1111110000001111",
    "1111110010101011",
    "1111111101100001",
    "1111110000111010",
    "1111011011010001",
    "1111000100001000",
    "1110101101111111",
    "1110011010111000",
    "1110001100100001",
    "1110000100000001",
    "1110000010000101",
    "1110000110110111",
    "1110010010001111",
    "1110100011101110",
    "1110111010100101",
    "1111010101011111",
    "1111110010100000",
    "1111110001000000",
    "1111010111111111",
    "1111000100111011",
    "1110111001010000",
    "1110110100101111",
    "1110110101101110",
    "1110111001011101",
    "1110111101010111",
    "1110111111110000",
    "1111000000011100",
    "1111000000011010",
    "1111000001010010",
    "1111000100011010",
    "1111001010010110",
    "1111010010101100",
    "1111011100001111",
    "1111100101100010",
    "1111101101001100",
    "1111110010011111",
    "1111110101011011",
    "1111110110101111",
    "1111110111101100",
    "1111111001110010",
    "1111111110010111",
    "1111111001100110",
    "1111101101111011",
    "1111011111000101",
    "1111001110010001",
    "1110111100111100",
    "1110101100101101",
    "1110011110111101",
    "1110010100100101",
    "1110001110001001",
    "1110001011101000",
    "1110001100111000",
    "1110010001011110",
    "1110011000101111",
    "1110100010001011",
    "1110101101010010",
    "1110111001110010",
    "1111000111101111",
    "1111010111010110",
    "1111101000111000",
    "1111111100001101",
    "1111101111010111",
    "1111011011011011",
    "1111001001111111",
    "1110111101000101",
    "1110110110001000",
    "1110110101100100",
    "1110111010110111",
    "1111000100111001",
    "1111010010010000",
    "1111100001011110",
    "1111110000111101",
    "1111111111000010",
    "1111110110000100",
    "1111110000001001",
    "1111110000100000",
    "1111110111111101",
    "1111111001101001",
    "1111100101110100",
    "1111001111001100",
    "1110111001000111",
    "1110100111000100",
    "1110011011110101",
    "1110011001000001",
    "1110011111000111",
    "1110101101011110",
    "1111000010110100",
    "1111011101000100",
    "1111111001001101",
    "1111101100000111",
    "1111010110011101",
    "1111001000010110",
    "1111000011000000",
    "1111000101111100",
    "1111001111101011",
    "1111011110001001",
    "1111101111101010",
    "1111111100111000",
    "1111101000011011",
    "1111010100000000",
    "1111000000111110",
    "1110110000111101",
    "1110100101011000",
    "1110011110111111",
    "1110011101100100",
    "1110011111111101",
    "1110100100011100",
    "1110101001100010",
    "1110101110101001",
    "1110110100000011",
    "1110111010101111",
    "1111000011101010",
    "1111001111011110",
    "1111011110000010",
    "1111101110110101",
    "1111111111000010",
    "1111101100110101",
    "1111011100000010",
    "1111001110001101",
    "1111000100110110",
    "1111000000110011",
    "1111000010000011",
    "1111000111101101",
    "1111010000010001",
    "1111011010000001",
    "1111100011101111",
    "1111101100111111",
    "1111110110000101",
    "1111111111111011",
    "1111110100101000",
    "1111100111011110",
    "1111011001011000",
    "1111001100000010",
    "1111000001100001",
    "1110111011010100",
    "1110111010000010",
    "1110111101000101",
    "1111000011000110",
    "1111001010100110",
    "1111010010100010",
    "1111011010101010",
    "1111100011000101",
    "1111101100000011",
    "1111110101010001",
    "1111111101110000",
    "1111111011110100",
    "1111111000111000",
    "1111111010000011",
    "1111111110111111",
    "1111111001101101",
    "1111110010001101",
    "1111101100101011",
    "1111101010110110",
    "1111101101100101",
    "1111110100101101",
    "1111111111001100",
    "1111110100100000",
    "1111101000001110",
    "1111011101011001",
    "1111010100111001",
    "1111001111000000",
    "1111001011011011",
    "1111001001011110",
    "1111001000100101",
    "1111001000011000",
    "1111001001000110",
    "1111001011011101",
    "1111010000101100",
    "1111011010001100",
    "1111101000101110",
    "1111111100001101",
    "1111101100101010",
    "1111010100011111",
    "1110111110011011",
    "1110101101100110",
    "1110100100001110",
    "1110100011000011",
    "1110101001010001",
    "1110110100111110",
    "1111000011100111",
    "1111010010110001",
    "1111100000100100",
    "1111101011111110",
    "1111110100100000",
    "1111111010001010",
    "1111111101000101",
    "1111111101100001",
    "1111111100000000",
    "1111111001001101",
    "1111110110000001",
    "1111110011010001",
    "1111110001011111",
    "1111110000110000",
    "1111110000110100",
    "1111110001001110",
    "1111110001101010",
    "1111110010000011",
    "1111110010110000",
    "1111110100100001",
    "1111111000001100",
    "1111111110010110",
    "1111111000111101",
    "1111101110100100",
    "1111100011110100",
    "1111011010011000",
    "1111010011101100",
    "1111010000110101",
    "1111010010001010",
    "1111010111100010",
    "1111100000100111",
    "1111101100111010",
    "1111111011111100",
    "1111110010110111",
    "1111100000100111",
    "1111001110111111",
    "1111000000001111",
    "1110110110111100",
    "1110110101011010",
    "1110111100111101",
    "1111001101001100",
    "1111100011111011",
    "1111111101011100",
    "1111101010100001",
    "1111010111111110",
    "1111001101100011",
    "1111001100010111",
    "1111010100001010",
    "1111100011101001",
    "1111111000111001",
    "1111101110100100",
    "1111010101101010",
    "1110111111010100",
    "1110101110000010",
    "1110100011011101",
    "1110100000000000",
    "1110100010110100",
    "1110101010001001",
    "1110110011111000",
    "1110111110001100",
    "1111000111101101",
    "1111001111101000",
    "1111010101011011",
    "1111011000110111",
    "1111011001111010",
    "1111011000110111",
    "1111010110011111",
    "1111010011110001",
    "1111010001111001",
    "1111010001111011",
    "1111010100011010",
    "1111011001011001",
    "1111100000110011",
    "1111101010011111",
    "1111110110100000",
    "1111111011001001",
    "1111101010111110",
    "1111011001111111",
    "1111001001100111",
    "1110111011010100",
    "1110110000010100",
    "1110101001001110",
    "1110100110000100",
    "1110100110101100",
    "1110101011000100",
    "1110110011101001",
    "1111000000111101",
    "1111010010111110",
    "1111101000100011",
    "1111111111001111",
    "1111101100000011",
    "1111011100010111",
    "1111010011100001",
    "1111010001101110",
    "1111010101101010",
    "1111011100111111",
    "1111100101011010",
    "1111101101001010",
    "1111110011011000",
    "1111110111101011",
    "1111111001111010",
    "1111111001111000",
    "1111110111011111",
    "1111110010110110",
    "1111101100011101",
    "1111100101001101",
    "1111011110001101",
    "1111011000100011",
    "1111010100111100",
    "1111010011101001",
    "1111010100011101",
    "1111010111001000",
    "1111011011100000",
    "1111100001100111",
    "1111101001110011",
    "1111110100001110",
    "1111111111001000",
    "1111110000111111",
    "1111100010011100",
    "1111010101000011",
    "1111001010011101",
    "1111000100000001",
    "1111000010110001",
    "1111000110111111",
    "1111010000011110",
    "1111011110010010",
    "1111101110111011",
    "1111111111101000",
    "1111101111101110",
    "1111100011011100",
    "1111011100010011",
    "1111011010110010",
    "1111011110010111",
    "1111100101011101",
    "1111101110000111",
    "1111110110100000",
    "1111111101011010",
    "1111111101101010",
    "1111111010101011",
    "1111111001001100",
    "1111111000110110",
    "1111111001011100",
    "1111111011000000",
    "1111111101100101",
    "1111111111000001",
    "1111111011010000",
    "1111110111101101",
    "1111110100111010",
    "1111110011001110",
    "1111110010101101",
    "1111110011010011",
    "1111110100110101",
    "1111110111001010",
    "1111111010001100",
    "1111111101110011",
    "1111111110000110",
    "1111111001101000",
    "1111110100100011",
    "1111101110100011",
    "1111100111011011",
    "1111011111011110",
    "1111010111101100",
    "1111010001100110",
    "1111001111000111",
    "1111010001110001",
    "1111011010001111",
    "1111100111110111",
    "1111111000101000",
    "1111110110010000",
    "1111100111110101",
    "1111011110011110",
    "1111011011011110",
    "1111011110111011",
    "1111100111111111",
    "1111110101001100",
    "1111111011000001",
    "1111101010001100",
    "1111011001101010",
    "1111001010110101",
    "1110111111001010",
    "1110110111110101",
    "1110110101100101",
    "1110111000010110",
    "1110111111000111",
    "1111000111111111",
    "1111010000110000",
    "1111010111001001",
    "1111011001100000",
    "1111010111001001",
    "1111010000011010",
    "1111000110101100",
    "1110111011110101",
    "1110110001111000",
    "1110101010100010",
    "1110100110111001",
    "1110100111010110",
    "1110101011101010",
    "1110110011000001",
    "1110111100100000",
    "1111000110110110",
    "1111010000110101",
    "1111011000111111",
    "1111011110000000",
    "1111011110100110",
    "1111011001111100",
    "1111010000001010",
    "1111000010001111",
    "1110110010000011",
    "1110100001111101",
    "1110010100000101",
    "1110001001111100",
    "1110000100000000",
    "1110000001101001",
    "1110000001100111",
    "1110000010100010",
    "1110000011011010",
    "1110000100100010",
    "1110001000000001",
    "1110010000111101",
    "1110100001100111",
    "1110111010000110",
    "1111010111100010",
    "1111110100110101",
    "1111110011101111",
    "1111100110110011",
    "1111100110000000",
    "1111101111110010",
    "1111111111011011",
    "1111101011110011",
    "1111011000101000",
    "1111000111111110",
    "1110111011000001",
    "1110110010101100",
    "1110110000000010",
    "1110110100011000",
    "1111000000111011",
    "1111010101100101",
    "1111110000100110",
    "1111110001011101",
    "1111010100111011",
    "1110111101100011",
    "1110101101100100",
    "1110100101010010",
    "1110100011010111",
    "1110100101101100",
    "1110101010001011",
    "1110101111011100",
    "1110110101001000",
    "1110111011110011",
    "1111000100100111",
    "1111010000100110",
    "1111011111111101",
    "1111110001111001",
    "1111111011011100",
    "1111101010100101",
    "1111011110000010",
    "1111010111101101",
    "1111011000011000",
    "1111011111100011",
    "1111101011101100",
    "1111111010011010",
    "1111110111000001",
    "1111101011011000",
    "1111100100100100",
    "1111100011011000",
    "1111100111100010",
    "1111101111110101",
    "1111111010110000",
    "1111111001001111",
    "1111101101101110",
    "1111100011111001",
    "1111011100110011",
    "1111011001001110",
    "1111011001011101",
    "1111011101010110",
    "1111100100000110",
    "1111101100010111",
    "1111110100100100",
    "1111111011010000",
    "1111111111100101",
    "1111111110010110",
    "1111111101110111",
    "1111111101110001",
    "1111111100111010",
    "1111111010101010",
    "1111110111000100",
    "1111110010111110",
    "1111101111101010",
    "1111101110100100",
    "1111110000111000",
    "1111110111001011",
    "1111111110110011",
    "1111110010010110",
    "1111100101010111",
    "1111011010000010",
    "1111010010011001",
    "1111001111110000",
    "1111010010101110",
    "1111011010111111",
    "1111100111101110",
    "1111110111101000",
    "1111110110101110",
    "1111100100111001",
    "1111010100100111",
    "1111000111110001",
    "1111000000001111",
    "1110111111011110",
    "1111000101111001",
    "1111010010100110",
    "1111100011001101",
    "1111110100011100",
    "1111111100111000",
    "1111110011001100",
    "1111101111011000",
    "1111110000110101",
    "1111110101111111",
    "1111111101000010",
    "1111111011011011",
    "1111110100010001",
    "1111101101101101",
    "1111100111110010",
    "1111100010101110",
    "1111011111000000",
    "1111011101010010",
    "1111011101111010",
    "1111100000101011",
    "1111100100101001",
    "1111101000100111",
    "1111101011001111",
    "1111101011100110",
    "1111101001011101",
    "1111100101001101",
    "1111011111110000",
    "1111011010010100",
    "1111010110001011",
    "1111010100010011",
    "1111010101010101",
    "1111011001001011",
    "1111011111000111",
    "1111100101111001",
    "1111101100000111",
    "1111110000011111",
    "1111110010010100",
    "1111110001011111",
    "1111101110011100",
    "1111101001110010",
    "1111100011111100",
    "1111011100110111",
    "1111010011111000",
    "1111001000001011",
    "1110111001000110",
    "1110100111000110",
    "1110010011111001",
    "1110000010001101",
    "1101110101000000",
    "1101101110100011",
    "1101110000000010",
    "1101111001010101",
    "1110001001100011",
    "1110011111101011",
    "1110111010011001",
    "1111010111111111",
    "1111110110000001",
    "1111101110101000",
    "1111011001001011",
    "1111001011110011",
    "1111000111011010",
    "1111001010111100",
    "1111010100000101",
    "1111100000001101",
    "1111101101011010",
    "1111111011000101",
    "1111110110010110",
    "1111100110011101",
    "1111010101010000",
    "1111000100000011",
    "1110110101000101",
    "1110101010110111",
    "1110100111001001",
    "1110101010000111",
    "1110110010011010",
    "1110111101101001",
    "1111001001001100",
    "1111010010110100",
    "1111011000111100",
    "1111011010101000",
    "1111010111100010",
    "1111001111110011",
    "1111000100000110",
    "1110110101100000",
    "1110100101011011",
    "1110010101100010",
    "1110000111100010",
    "1101111100110010",
    "1101110110001011",
    "1101110011110100",
    "1101110101001110",
    "1101111001101111",
    "1110000000100100",
    "1110001001100101",
    "1110010101011101",
    "1110100101000101",
    "1110111000101111",
    "1111001111011110",
    "1111100110101011",
    "1111111010111011",
    "1111110111001100",
    "1111110010000100",
    "1111110110001000",
    "1111111110001010",
    "1111101101101101",
    "1111011011101111",
    "1111001010111000",
    "1110111100110010",
    "1110110001111110",
    "1110101010011000",
    "1110100101101001",
    "1110100011100010",
    "1110100011111110",
    "1110100110110111",
    "1110101100001010",
    "1110110011110100",
    "1110111101111111",
    "1111001010111101",
    "1111011011001001",
    "1111101110101000",
    "1111111011001010",
    "1111100100000101",
    "1111001110101001",
    "1110111101100011",
    "1110110010100010",
    "1110101110000000",
    "1110101111000010",
    "1110110011110100",
    "1110111010100011",
    "1111000010000110",
    "1111001010001001",
    "1111010010100100",
    "1111011010110101",
    "1111100001011010",
    "1111100011111011",
    "1111100000000011",
    "1111010100100100",
    "1111000010001101",
    "1110101011110010",
    "1110010101011000",
    "1110000011001101",
    "1101111000010110",
    "1101110110010011",
    "1101111100111010",
    "1110001011001111",
    "1110100000000000",
    "1110111001100101",
    "1111010101111001",
    "1111110010001101",
    "1111110100101101",
    "1111100001110011",
    "1111010110110110",
    "1111010011101110",
    "1111010110100101",
    "1111011100011011",
    "1111100010001011",
    "1111100101111011",
    "1111100111010000",
    "1111100111001100",
    "1111100111011001",
    "1111101001100001",
    "1111101110011010",
    "1111110110001011",
    "1111111111100011",
    "1111110011011100",
    "1111100101101110",
    "1111010110011111",
    "1111000101111001",
    "1110110100100000",
    "1110100011100110",
    "1110010100110011",
    "1110001001101010",
    "1110000010111101",
    "1110000000011111",
    "1110000001001101",
    "1110000011100111",
    "1110000110011000",
    "1110001000110000",
    "1110001010111000",
    "1110001101100011",
    "1110010001101100",
    "1110011000001011",
    "1110100001001111",
    "1110101100011100",
    "1110111000111001",
    "1111000101001001",
    "1111001111111000",
    "1111010111111100",
    "1111011100101110",
    "1111011110001111",
    "1111011101001010",
    "1111011010110111",
    "1111011000111111",
    "1111011001011000",
    "1111011101001111",
    "1111100101001001",
    "1111110000011010",
    "1111111101011101",
    "1111110101110000",
    "1111101011011010",
    "1111100101000011",
    "1111100011100100",
    "1111100111001110",
    "1111101111100111",
    "1111111100000011",
    "1111110100100000",
    "1111100011110100",
    "1111010011111011",
    "1111000111001110",
    "1110111111110011",
    "1110111111000111",
    "1111000101100100",
    "1111010010100010",
    "1111100100011100",
    "1111111000111010",
    "1111110010100001",
    "1111100000001100",
    "1111010001100001",
    "1111000111000100",
    "1111000000011100",
    "1110111100100101",
    "1110111010001111",
    "1110111000100000",
    "1110110111001110",
    "1110110111000100",
    "1110111001010110",
    "1110111111011010",
    "1111001010000010",
    "1111011001000001",
    "1111101010111101",
    "1111111101100110",
    "1111110001101010",
    "1111100101001101",
    "1111011110010110",
    "1111011101010010",
    "1111100001000101",
    "1111100111111101",
    "1111101111101110",
    "1111110110010000",
    "1111111001110010",
    "1111111001001110",
    "1111110100010000",
    "1111101011010001",
    "1111011111010111",
    "1111010010000011",
    "1111000101000101",
    "1110111010000100",
    "1110110010010000",
    "1110101110010001",
    "1110101101111010",
    "1110110000010111",
    "1110110100100000",
    "1110111001001110",
    "1110111101101110",
    "1111000001101100",
    "1111000101001110",
    "1111001000101111",
    "1111001100110000",
    "1111010001111000",
    "1111011000110101",
    "1111100010010101",
    "1111101110111111",
    "1111111110111011",
    "1111101110100110",
    "1111011011011110",
    "1111001010100010",
    "1110111110111010",
    "1110111011010100",
    "1111000001001100",
    "1111010000010010",
    "1111100110110011",
    "1111111110010010",
    "1111100010110011",
    "1111001010010001",
    "1110110111100010",
    "1110101100001010",
    "1110101000101000",
    "1110101100001001",
    "1110110101010010",
    "1111000010010010",
    "1111010001100010",
    "1111100001100001",
    "1111110001000010",
    "1111111110111111",
    "1111110101011000",
    "1111101100011100",
    "1111100110000000",
    "1111100001010111",
    "1111011101101000",
    "1111011001111100",
    "1111010101101100",
    "1111010000101100",
    "1111001011010011",
    "1111000101111110",
    "1111000001011110",
    "1110111110010110",
    "1110111101000000",
    "1110111101101011",
    "1111000000010111",
    "1111000101000101",
    "1111001011110011",
    "1111010100011100",
    "1111011110110101",
    "1111101010110000",
    "1111110111111001",
    "1111111010000110",
    "1111101011111001",
    "1111011110001111",
    "1111010001111110",
    "1111000111111110",
    "1111000000110110",
    "1110111101000000",
    "1110111100011110",
    "1110111111000100",
    "1111000100011010",
    "1111001100001001",
    "1111010101101001",
    "1111011111111111",
    "1111101010000000",
    "1111110010010011",
    "1111110111100000",
    "1111111000100111",
    "1111110101010100",
    "1111101110010010",
    "1111100101001101",
    "1111011100100000",
    "1111010110101010",
    "1111010101110100",
    "1111011011000100",
    "1111100110100100",
    "1111110111011100",
    "1111110011111001",
    "1111011101101101",
    "1111001000011000",
    "1110110110001000",
    "1110101000101000",
    "1110100000101100",
    "1110011110001100",
    "1110100000001000",
    "1110100101001000",
    "1110101011110010",
    "1110110011001101",
    "1110111011001010",
    "1111000100000011",
    "1111001110100100",
    "1111011011011110",
    "1111101011000001",
    "1111111100101100",
    "1111110000110011",
    "1111011111011111",
    "1111010001010010",
    "1111000111101010",
    "1111000011010000",
    "1111000011111000",
    "1111001000011101",
    "1111001111100100",
    "1111010111100111",
    "1111011111001101",
    "1111100101010101",
    "1111101001100001",
    "1111101011110011",
    "1111101100100110",
    "1111101100101010",
    "1111101100111100",
    "1111101110010111",
    "1111110001110000",
    "1111110111101000",
    "1111111111111101",
    "1111110101110110",
    "1111101011000111",
    "1111100001010100",
    "1111011001110100",
    "1111010101011000",
    "1111010100001010",
    "1111010101011111",
    "1111011000010011",
    "1111011011100001",
    "1111011110010110",
    "1111100000010100",
    "1111100001010111",
    "1111100001110001",
    "1111100001111101",
    "1111100010010101",
    "1111100011011101",
    "1111100101111011",
    "1111101010011000",
    "1111110001100011",
    "1111111011111100",
    "1111110110011110",
    "1111100110110100",
    "1111010111001000",
    "1111001010000100",
    "1111000010001010",
    "1111000000111101",
    "1111000110101000",
    "1111010010000000",
    "1111100000111110",
    "1111110001001101",
    "1111111111001010",
    "1111110001100010",
    "1111100110110000",
    "1111011111011111",
    "1111011100011100",
    "1111011110000101",
    "1111100100010010",
    "1111101110000001",
    "1111111001011010",
    "1111111011110101",
    "1111110100000001",
    "1111110000100101",
    "1111110001111101",
    "1111110111100111",
    "1111111111100110",
    "1111110101000011",
    "1111101001111001",
    "1111011111010010",
    "1111010110010010",
    "1111010000000010",
    "1111001101011100",
    "1111001111000100",
    "1111010100110100",
    "1111011110000000",
    "1111101001010010",
    "1111110101000101",
    "1111111111111101",
    "1111110111000101",
    "1111110000101011",
    "1111101100110101",
    "1111101011011011",
    "1111101100000111",
    "1111101110100010",
    "1111110010010000",
    "1111110110101101",
    "1111111011010001",
    "1111111111010000",
    "1111111101110011",
    "1111111100001111",
    "1111111011111010",
    "1111111100010111",
    "1111111101000110",
    "1111111101100111",
    "1111111101100101",
    "1111111100110010",
    "1111111011000001",
    "1111111000000001",
    "1111110011011101",
    "1111101101001001",
    "1111100101011000",
    "1111011100111100",
    "1111010101001101",
    "1111001111110000",
    "1111001101111101",
    "1111010000101011",
    "1111011000010001",
    "1111100100101110",
    "1111110101011110",
    "1111110110100001",
    "1111100001001111",
    "1111001100111111",
    "1110111100010001",
    "1110110001000101",
    "1110101100011011",
    "1110101101111011",
    "1110110100001010",
    "1110111100111111",
    "1111000110011111",
    "1111001111100100",
    "1111011000011101",
    "1111100010000101",
    "1111101101101101",
    "1111111011110101",
    "1111110100000011",
    "1111100011101001",
    "1111010101000001",
    "1111001010001011",
    "1111000100000110",
    "1111000010101111",
    "1111000101001101",
    "1111001001111111",
    "1111001111101011",
    "1111010101000001",
    "1111011001001011",
    "1111011011100000",
    "1111011011101101",
    "1111011001100111",
    "1111010101000011",
    "1111001101111111",
    "1111000100101100",
    "1110111001111010",
    "1110101110110011",
    "1110100100110110",
    "1110011101010111",
    "1110011001011001",
    "1110011001011001",
    "1110011101010010",
    "1110100100100101",
    "1110101110100100",
    "1110111010011110",
    "1111000111100011",
    "1111010101001001",
    "1111100010101110",
    "1111101111110011",
    "1111111011111011",
    "1111111001010010",
    "1111110000010100",
    "1111101001100010",
    "1111100101010000",
    "1111100011101010",
    "1111100100111011",
    "1111101001000101",
    "1111110000000111",
    "1111111001111100",
    "1111111001101001",
    "1111101011011101",
    "1111011100101010",
    "1111001111000100",
    "1111000100111001",
    "1111000000010001",
    "1111000010101011",
    "1111001100101101",
    "1111011101101001",
    "1111110011100001",
    "1111110100100100",
    "1111011110001001",
    "1111001100001111",
    "1111000001000101",
    "1110111101100110",
    "1111000001100111",
    "1111001100011100",
    "1111011101010001",
    "1111110011000110",
    "1111110011110000",
    "1111011001111010",
    "1111000010011001",
    "1110110000000101",
    "1110100100111001",
    "1110100001000101",
    "1110100011010011",
    "1110101001000111",
    "1110110000001010",
    "1110110111000011",
    "1110111101011100",
    "1111000011101001",
    "1111001001111001",
    "1111001111110011",
    "1111010100001011",
    "1111010101011101",
    "1111010010010111",
    "1111001010101101",
    "1110111111100110",
    "1110110011001111",
    "1110101000000001",
    "1110011111110110",
    "1110011011100011",
    "1110011011000100",
    "1110011101101101",
    "1110100010110011",
    "1110101001101111",
    "1110110010000101",
    "1110111011100001",
    "1111000101110110",
    "1111010000110011",
    "1111011100001111",
    "1111101000001011",
    "1111110100110100",
    "1111111101001101",
    "1111101101010010",
    "1111011011000010",
    "1111000110111111",
    "1110110010101011",
    "1110100000001010",
    "1110010001100100",
    "1110001000001110",
    "1110000100011100",
    "1110000101010011",
    "1110001001001011",
    "1110001110001111",
    "1110010011001000",
    "1110010111000110",
    "1110011010101011",
    "1110100000001100",
    "1110101010110000",
    "1110111100100001",
    "1111010101010000",
    "1111110001100110",
    "1111110011101101",
    "1111100000001010",
    "1111010111100011",
    "1111011010011001",
    "1111100101111011",
    "1111110101011011",
    "1111111011101001",
    "1111110000011110",
    "1111101001111110",
    "1111100111100010",
    "1111100111110110",
    "1111101001110001",
    "1111101100111010",
    "1111110001011101",
    "1111110111100100",
    "1111111111000001",
    "1111111001001010",
    "1111110010011011",
    "1111101101111111",
    "1111101100010000",
    "1111101100110011",
    "1111101110101101",
    "1111110001000110",
    "1111110011100010",
    "1111110101111111",
    "1111111000111000",
    "1111111100110100",
    "1111111101110010",
    "1111110111000011",
    "1111101111100010",
    "1111101000010101",
    "1111100010101011",
    "1111011111100110",
    "1111011111110001",
    "1111100011010000",
    "1111101001100001",
    "1111110001100111",
    "1111111010001101",
    "1111111110001100",
    "1111111001010101",
    "1111111000110110",
    "1111111110000101",
    "1111110110010001",
    "1111100100100111",
    "1111001110011001",
    "1110110101110111",
    "1110011101100110",
    "1110000111111110",
    "1101110110101100",
    "1101101010100101",
    "1101100011101100",
    "1101100001010100",
    "1101100010100010",
    "1101100110010110",
    "1101101011111000",
    "1101110010010101",
    "1101111001011000",
    "1110000001000011",
    "1110001001110010",
    "1110010011111000",
    "1110011111001101",
    "1110101011000100",
    "1110110110000100",
    "1110111110100001",
    "1111000010101111",
    "1111000001101011",
    "1110111011000111",
    "1110110000000010",
    "1110100010010100",
    "1110010100011010",
    "1110001000110000",
    "1110000001010010",
    "1101111111000100",
    "1110000010011001",
    "1110001011001001",
    "1110011001011000",
    "1110101101011100",
    "1111000111101000",
    "1111100110111111",
    "1111110111010010",
    "1111010111101100",
    "1110111111000000",
    "1110110001000010",
    "1110101111001100",
    "1110111000000100",
    "1111001000010110",
    "1111011100010100",
    "1111110001010111",
    "1111111001010101",
    "1111100011101010",
    "1111001101110010",
    "1110111000111100",
    "1110100111110001",
    "1110011101011001",
    "1110011100010100",
    "1110100101011011",
    "1110110111101101",
    "1111010000010101",
    "1111101011101111",
    "1111111001100111",
    "1111100010100001",
    "1111010000101110",
    "1111000100111001",
    "1110111111000111",
    "1110111110101110",
    "1111000010101001",
    "1111001001011001",
    "1111010001011110",
    "1111011001011001",
    "1111100000001100",
    "1111100101010010",
    "1111101000101010",
    "1111101010101100",
    "1111101011111010",
    "1111101100110110",
    "1111101101111110",
    "1111101111110001",
    "1111110010110111",
    "1111110111110101",
    "1111111110111010",
    "1111111000010010",
    "1111101110110010",
    "1111100110000001",
    "1111011111011001",
    "1111011011110111",
    "1111011011100101",
    "1111011110000010",
    "1111100010010000",
    "1111100111100110",
    "1111101101111111",
    "1111110101110110",
    "1111111111110100",
    "1111110011111000",
    "1111100110000100",
    "1111011000011011",
    "1111001101011001",
    "1111000111010101",
    "1111000111110100",
    "1111001111001100",
    "1111011100001110",
    "1111101100100011",
    "1111111101011000",
    "1111110011110110",
    "1111101001000000",
    "1111100010111001",
    "1111100001011111",
    "1111100100001010",
    "1111101010001011",
    "1111110010110110",
    "1111111101100000",
    "1111110110101101",
    "1111101011010000",
    "1111100001111011",
    "1111011100101011",
    "1111011100111111",
    "1111100011001010",
    "1111101110001101",
    "1111111100000000",
    "1111110110001101",
    "1111101010111000",
    "1111100011011100",
    "1111100000000111",
    "1111100000000111",
    "1111100010010101",
    "1111100101111110",
    "1111101010101111",
    "1111110001000101",
    "1111111001111001",
    "1111111001111111",
    "1111101010011001",
    "1111011000000011",
    "1111000100110011",
    "1110110011001010",
    "1110100101101111",
    "1110011110110001",
    "1110011111010100",
    "1110100111001101",
    "1110110100111100",
    "1111000110001110",
    "1111011000011101",
    "1111101001010011",
    "1111110111000011",
    "1111111111010011",
    "1111111010001010",
    "1111111001010101",
    "1111111100001100",
    "1111111110000101",
    "1111110110100111",
    "1111101110100001",
    "1111100110111000",
    "1111100000100100",
    "1111011100001001",
    "1111011001110010",
    "1111011001001110",
    "1111011001111101",
    "1111011011011101",
    "1111011101001100",
    "1111011110111111",
    "1111100000111001",
    "1111100011011100",
    "1111100111000111",
    "1111101100011000",
    "1111110011001000",
    "1111111010100001",
    "1111111110110100",
    "1111111010101011",
    "1111111010100000",
    "1111111111001101",
    "1111110111001000",
    "1111101001010101",
    "1111011000101000",
    "1111000110011000",
    "1110110011111011",
    "1110100010100111",
    "1110010100000001",
    "1110001010000001",
    "1110000110110001",
    "1110001100000010",
    "1110011010101011",
    "1110110001110000",
    "1111001110011111",
    "1111101100101110",
    "1111110111111110",
    "1111100011001111",
    "1111010110110111",
    "1111010010101111",
    "1111010101010011",
    "1111011100011100",
    "1111100110011110",
    "1111110010011101",
    "1111111111110011",
    "1111110000100101",
    "1111100000011110",
    "1111010000110001",
    "1111000011011010",
    "1110111010001110",
    "1110110110011000",
    "1110110111111001",
    "1110111101011110",
    "1111000101000000",
    "1111001011111010",
    "1111010000000010",
    "1111010000000000",
    "1111001011100001",
    "1111000011010011",
    "1110111000101101",
    "1110101101010001",
    "1110100010100010",
    "1110011001100111",
    "1110010011001010",
    "1110001111011001",
    "1110001110010001",
    "1110001111011111",
    "1110010010111101",
    "1110011000110010",
    "1110100001101001",
    "1110101110010100",
    "1110111111001010",
    "1111010011100110",
    "1111101001111100",
    "1111111111100110",
    "1111101110010000",
    "1111100010001000",
    "1111011101010010",
    "1111011111101100",
    "1111100111111110",
    "1111110011111001",
    "1111111111000100",
    "1111110011010110",
    "1111101010110110",
    "1111100110110000",
    "1111100111100111",
    "1111101101001111",
    "1111110110101100",
    "1111111101101101",
    "1111110010010111",
    "1111101001110110",
    "1111100110011101",
    "1111101001101101",
    "1111110011111101",
    "1111111011110011",
    "1111100111111011",
    "1111010011010000",
    "1111000000101100",
    "1110110010100010",
    "1110101010000100",
    "1110100111011000",
    "1110101001101010",
    "1110101111100100",
    "1110110111111001",
    "1111000001100111",
    "1111001100001111",
    "1111010111011011",
    "1111100010110110",
    "1111101101111011",
    "1111110111111100",
    "1111111111111011",
    "1111111010010111",
    "1111110111101010",
    "1111110111101011",
    "1111111001111011",
    "1111111101101100",
    "1111111101110000",
    "1111111001001011",
    "1111110101001011",
    "1111110010011111",
    "1111110001111111",
    "1111110100110011",
    "1111111011111001",
    "1111111000001100",
    "1111100111111111",
    "1111010100111011",
    "1111000001010010",
    "1110101111100011",
    "1110100001101110",
    "1110011001000100",
    "1110010101101100",
    "1110010110110111",
    "1110011011010110",
    "1110100001101110",
    "1110101000110101",
    "1110101111101100",
    "1110110101101001",
    "1110111010000110",
    "1110111100110101",
    "1110111101110111",
    "1110111101011110",
    "1110111100011001",
    "1110111011011001",
    "1110111011001100",
    "1110111100001001",
    "1110111101111111",
    "1111000000000000",
    "1111000001000000",
    "1110111111111000",
    "1110111011101111",
    "1110110100001110",
    "1110101001110100",
    "1110011101101101",
    "1110010001110011",
    "1110001000010101",
    "1110000011001101",
    "1110000011101010",
    "1110001001111101",
    "1110010101011011",
    "1110100100110001",
    "1110110110011111",
    "1111001001001011",
    "1111011011100101",
    "1111101100100111",
    "1111111011001010",
    "1111111001110010",
    "1111110011000110",
    "1111110000111101",
    "1111110010110110",
    "1111110111010111",
    "1111111100011111",
    "1111111111111101",
    "1111111111111000",
    "1111111011010001",
    "1111110010011010",
    "1111100110110010",
    "1111011010100101",
    "1111010000001000",
    "1111001001010000",
    "1111000110111110",
    "1111001001010110",
    "1111001111110000",
    "1111011001001110",
    "1111100100101110",
    "1111110001011101",
    "1111111110110100",
    "1111110011110001",
    "1111100111001111",
    "1111011100101110",
    "1111010101011111",
    "1111010010101111",
    "1111010101001000",
    "1111011100010111",
    "1111100111010111",
    "1111110100000111",
    "1111111111100000",
    "1111110101100101",
    "1111101111100001",
    "1111101101111011",
    "1111110000101010",
    "1111110111000000",
    "1111111111110001",
    "1111110110011000",
    "1111101101000010",
    "1111100101101010",
    "1111100001110110",
    "1111100010111001",
    "1111101001101001",
    "1111110101111111",
    "1111111001011011",
    "1111100110111101",
    "1111010101011000",
    "1111000111010001",
    "1110111110011011",
    "1110111011011000",
    "1110111101011100",
    "1111000011000000",
    "1111001010001100",
    "1111010001100001",
    "1111011000011011",
    "1111100000000101",
    "1111101010111101",
    "1111111011010101",
    "1111101110000101",
    "1111010011010101",
    "1110111000101000",
    "1110100011010010",
    "1110010111111110",
    "1110011001010001",
    "1110100110111100",
    "1110111110001100",
    "1111011010110000",
    "1111110111111000",
    "1111101110010101",
    "1111011010101101",
    "1111001110010111",
    "1111001001000110",
    "1111001001110010",
    "1111001110111010",
    "1111010110110111",
    "1111100000100011",
    "1111101011000010",
    "1111110101101011",
    "1111111111110011",
    "1111110111001000",
    "1111101111101011",
    "1111101010000110",
    "1111100110100110",
    "1111100101000110",
    "1111100101001000",
    "1111100110000001",
    "1111100110111010",
    "1111100111000100",
    "1111100110000100",
    "1111100011101110",
    "1111011111111000",
    "1111011010100000",
    "1111010011100010",
    "1111001011000110",
    "1111000001011010",
    "1110110110111111",
    "1110101100011100",
    "1110100010101011",
    "1110011010100011",
    "1110010101001011",
    "1110010011010101",
    "1110010101100000",
    "1110011011101011",
    "1110100101011010",
    "1110110010000011",
    "1111000000111110",
    "1111010001110000",
    "1111100100000011",
    "1111110111011010",
    "1111110100111111",
    "1111100010101011",
    "1111010011001000",
    "1111000111110100",
    "1111000001100001",
    "1111000000000101",
    "1111000010100010",
    "1111000111011000",
    "1111001101001110",
    "1111010011011100",
    "1111011010010011",
    "1111100010100111",
    "1111101101011101",
    "1111111011001111",
    "1111110100101010",
    "1111100100001010",
    "1111010101111100",
    "1111001100111000",
    "1111001011000111",
    "1111010001011111",
    "1111011111001000",
    "1111110001100101",
    "1111111010101100",
    "1111101001100001",
    "1111011110000101",
    "1111011010100101",
    "1111011111111111",
    "1111101101111010",
    "1111111101010110",
    "1111100100111110",
    "1111001100110111",
    "1110111000111001",
    "1110101100001100",
    "1110101000010110",
    "1110101101010001",
    "1110111001010000",
    "1111001010000001",
    "1111011101100100",
    "1111110010110100",
    "1111110110100101",
    "1111011110110101",
    "1111000110100111",
    "1110101111101001",
    "1110011100010001",
    "1110001110101011",
    "1110001000000001",
    "1110000111111110",
    "1110001100110111",
    "1110010100001110",
    "1110011011111101",
    "1110100011000011",
    "1110101001101111",
    "1110110001010100",
    "1110111011011001",
    "1111001001100011",
    "1111011100100000",
    "1111110011110011",
    "1111110010001101",
    "1111011000100000",
    "1111000010010101",
    "1110110010100001",
    "1110101010011110",
    "1110101010000010",
    "1110101111100100",
    "1110111000100101",
    "1111000010110011",
    "1111001100111000",
    "1111010110111110",
    "1111100010011100",
    "1111110000111000",
    "1111111100110101",
    "1111100111101010",
    "1111010010000011",
    "1110111111010110",
    "1110110010100001",
    "1110101101000100",
    "1110101110110001",
    "1110110110001000",
    "1111000001010100",
    "1111001111001101",
    "1111011111011110",
    "1111110010000010",
    "1111111001110010",
    "1111100101111110",
    "1111010101010011",
    "1111001010110000",
    "1111001000100000",
    "1111001111000101",
    "1111011101001010",
    "1111101111110101",
    "1111111100011111",
    "1111101011100000",
    "1111100000000111",
    "1111011100000111",
    "1111100000010111",
    "1111101100011000",
    "1111111110100001",
    "1111101011111100",
    "1111010110011011",
    "1111000100001000",
    "1110110111010101",
    "1110110000111000",
    "1110110000010001",
    "1110110011111011",
    "1110111010000111",
    "1111000001101110",
    "1111001010011110",
    "1111010100111110",
    "1111100010000110",
    "1111110010011001",
    "1111111010011001",
    "1111100101011111",
    "1111010000101110",
    "1110111110010010",
    "1110110000001100",
    "1110100111110010",
    "1110100101101110",
    "1110101001110000",
    "1110110011000000",
    "1111000000000011",
    "1111001111010001",
    "1111011110110000",
    "1111101100111011",
    "1111111000011101",
    "1111111111001111",
    "1111111010001010",
    "1111110111101010",
    "1111110110110000",
    "1111110110100000",
    "1111110110010100",
    "1111110110000000",
    "1111110101101010",
    "1111110101011100",
    "1111110101011001",
    "1111110101010101",
    "1111110101000110",
    "1111110100100101",
    "1111110011110111",
    "1111110011000010",
    "1111110010000110",
    "1111110000110101",
    "1111101110110011",
    "1111101011100111",
    "1111100111001110",
    "1111100010000101",
    "1111011101000100",
    "1111011001010101",
    "1111010111111010",
    "1111011001011110",
    "1111011110001111",
    "1111100110000110",
    "1111110001001100",
    "1111111111111010",
    "1111101100101010",
    "1111010101001110",
    "1110111011100001",
    "1110100011000011",
    "1110010000000111",
    "1110000110010011",
    "1110000111011010",
    "1110010010111001",
    "1110100110011011",
    "1110111110111000",
    "1111011001010101",
    "1111110011100110",
    "1111110100000111",
    "1111011111110000",
    "1111010001001010",
    "1111001010000001",
    "1111001011000110",
    "1111010011110110",
    "1111100010101001",
    "1111110100111010",
    "1111110111110001",
    "1111100101010011",
    "1111010100100101",
    "1111000101110100",
    "1110111000111001",
    "1110101101110101",
    "1110100101000000",
    "1110011110110001",
    "1110011011010110",
    "1110011010010011",
    "1110011010110010",
    "1110011011111100",
    "1110011101010001",
    "1110011110110011",
    "1110100001000010",
    "1110100100100101",
    "1110101001110101",
    "1110110000110001",
    "1110111001000110",
    "1111000010011010",
    "1111001100100011",
    "1111010111011011",
    "1111100011000110",
    "1111101111011001",
    "1111111011101101",
    "1111111000111010",
    "1111101111101001",
    "1111101001010100",
    "1111100110000100",
    "1111100101010111",
    "1111100110000000",
    "1111100110110001",
    "1111100110110101",
    "1111100110000001",
    "1111100100101001",
    "1111100011001101",
    "1111100010000000",
    "1111100000111001",
    "1111011111011110",
    "1111011101000100",
    "1111011001011101",
    "1111010100110100",
    "1111010000000000",
    "1111001100001111",
    "1111001010110111",
    "1111001100111101",
    "1111010011010000",
    "1111011110000111",
    "1111101101011011",
    "1111111111010110",
    "1111101001100010",
    "1111010011001000",
    "1110111110110101",
    "1110101111011100",
    "1110100111010101",
    "1110100111100101",
    "1110101111110000",
    "1110111101111011",
    "1111001111010010",
    "1111100000101110",
    "1111101111100101",
    "1111111010001001",
    "1111111111101000",
    "1111111111110011",
    "1111111100011101",
    "1111110101101010",
    "1111101100111111",
    "1111100011100100",
    "1111011010001110",
    "1111010001011111",
    "1111001001101010",
    "1111000010110110",
    "1110111101000100",
    "1110111000010001",
    "1110110100100101",
    "1110110010010010",
    "1110110010000000",
    "1110110100100100",
    "1110111010101111",
    "1111000100101111",
    "1111010010010000",
    "1111100010000010",
    "1111110010010000",
    "1111111111000001",
    "1111110011101000",
    "1111101100101000",
    "1111101010001101",
    "1111101011110011",
    "1111110000010100",
    "1111110110100000",
    "1111111101001100",
    "1111111100011101",
    "1111110111000101",
    "1111110010111101",
    "1111110000010011",
    "1111101111010111",
    "1111110000011000",
    "1111110011100100",
    "1111111001001010",
    "1111111110101101",
    "1111110011111010",
    "1111100110000110",
    "1111010101000001",
    "1111000000111110",
    "1110101011001110",
    "1110010101110110",
    "1110000011011111",
    "1101110110110100",
    "1101110001100110",
    "1101110100010000",
    "1101111101101011",
    "1110001011101000",
    "1110011100010110",
    "1110110000000101",
    "1111001000011011",
    "1111100110011000",
    "1111110111001110",
    "1111010100011101",
    "1110110111000110",
    "1110100100101001",
    "1110100000011001",
    "1110101001101010",
    "1110111011111101",
    "1111010001000011",
    "1111100011010011",
    "1111101111101111",
    "1111110110001111",
    "1111111000010110",
    "1111111000001000",
    "1111110111000001",
    "1111110101010000",
    "1111110010011000",
    "1111101101111001",
    "1111101000000101",
    "1111100010001000",
    "1111011101110111",
    "1111011100110010",
    "1111011111010111",
    "1111100101000110",
    "1111101100111110",
    "1111110110000101",
    "1111111111101100",
    "1111110110101111",
    "1111101101111001",
    "1111100110011001",
    "1111100000110001",
    "1111011101010110",
    "1111011100000100",
    "1111011100011100",
    "1111011101101110",
    "1111011111000101",
    "1111011111111111",
    "1111100000001111",
    "1111011111110101",
    "1111011110101101",
    "1111011100100001",
    "1111011000110000",
    "1111010010111101",
    "1111001010111010",
    "1111000001001101",
    "1110110111001001",
    "1110101110011100",
    "1110101000100101",
    "1110100110010011",
    "1110100111100011",
    "1110101011110011",
    "1110110010011101",
    "1110111011000010",
    "1111000100111001",
    "1111001111001101",
    "1111011000110010",
    "1111100000000101",
    "1111100011011000",
    "1111100001001101",
    "1111011000110101",
    "1111001010111000",
    "1110111001010101",
    "1110100110111001",
    "1110010110011000",
    "1110001001111111",
    "1110000010111011",
    "1110000001001101",
    "1110000011110110",
    "1110001001011000",
    "1110010000011111",
    "1110011000001011",
    "1110011111110101",
    "1110100111010000",
    "1110101110010111",
    "1110110101001000",
    "1110111011011001",
    "1111000000111101",
    "1111000101011111",
    "1111001000110111",
    "1111001011001100",
    "1111001100110101",
    "1111001110001111",
    "1111001111111010",
    "1111010010001011",
    "1111010101011011",
    "1111011001111001",
    "1111011111110110",
    "1111100111011001",
    "1111110000011111",
    "1111111010101100",
    "1111111010101000",
    "1111110000011100",
    "1111100111101010",
    "1111100001000000",
    "1111011100111101",
    "1111011011101000",
    "1111011100110000",
    "1111011111110110",
    "1111100100001101",
    "1111101001001011",
    "1111101110001001",
    "1111110010101010",
    "1111110110100010",
    "1111111001110010",
    "1111111100100011",
    "1111111111000100",
    "1111111110011011",
    "1111111011111010",
    "1111111001011101",
    "1111110111100000",
    "1111110110101011",
    "1111110111110101",
    "1111111011110000",
    "1111111101000000",
    "1111110010101010",
    "1111100110001011",
    "1111011001010000",
    "1111001101110111",
    "1111000101110010",
    "1111000010000110",
    "1111000010111011",
    "1111000111100101",
    "1111001111000101",
    "1111011000101101",
    "1111100100010010",
    "1111110001111001",
    "1111111110011001",
    "1111101101011011",
    "1111011101000101",
    "1111010000000000",
    "1111001000111001",
    "1111001001100000",
    "1111010010001010",
    "1111100001011100",
    "1111110100110001",
    "1111110111000101",
    "1111100101011000",
    "1111011000110000",
    "1111010011000000",
    "1111010100111110",
    "1111011110010110",
    "1111101101100101",
    "1111111111110110",
    "1111101101001101",
    "1111011101011110",
    "1111010010111000",
    "1111001110011100",
    "1111001111111111",
    "1111010110011011",
    "1111100000011111",
    "1111101100111110",
    "1111111010111101",
    "1111110110010101",
    "1111100111111101",
    "1111011011001110",
    "1111010001101011",
    "1111001100101110",
    "1111001101001001",
    "1111010010100110",
    "1111011011101011",
    "1111100110010000",
    "1111110000000101",
    "1111110111010110",
    "1111111011001000",
    "1111111011100000",
    "1111111001011100",
    "1111110110010100",
    "1111110011101101",
    "1111110010111111",
    "1111110101000110",
    "1111111010011001",
    "1111111101010010",
    "1111110010111111",
    "1111100111111111",
    "1111011101110111",
    "1111010101111100",
    "1111010001000101",
    "1111001111011110",
    "1111010000101011",
    "1111010100000011",
    "1111011001000001",
    "1111011111011001",
    "1111100111011101",
    "1111110001111001",
    "1111111111000110",
    "1111110001010010",
    "1111100000110001",
    "1111010001100010",
    "1111000110000011",
    "1111000000010101",
    "1111000001110001",
    "1111001010101111",
    "1111011010100010",
    "1111101111010010",
    "1111111001111000",
    "1111100100100000",
    "1111010011101110",
    "1111001001110000",
    "1111000111001101",
    "1111001011000001",
    "1111010011000101",
    "1111011101001110",
    "1111101000001111",
    "1111110100010100",
    "1111111101100110",
    "1111101100110001",
    "1111011001011001",
    "1111000101000101",
    "1110110010100111",
    "1110100101001011",
    "1110011111010001",
    "1110100001110000",
    "1110101011110000",
    "1110111010111000",
    "1111001100000001",
    "1111011100001110",
    "1111101001010110",
    "1111110010010010",
    "1111110110110010",
    "1111110111001110",
    "1111110100010110",
    "1111101110101110",
    "1111100110100010",
    "1111011011101010",
    "1111001101110011",
    "1110111101001100",
    "1110101010111010",
    "1110011000110111",
    "1110001001100000",
    "1101111111010010",
    "1101111011110101",
    "1101111111101110",
    "1110001010001111",
    "1110011001110101",
    "1110101100100101",
    "1111000000110101",
    "1111010101010011",
    "1111101001001101",
    "1111111011111010",
    "1111110011001111",
    "1111100101010000",
    "1111011011001100",
    "1111010101111001",
    "1111010101101111",
    "1111011010010110",
    "1111100010110001",
    "1111101101110010",
    "1111111010100000",
    "1111110111011001",
    "1111101000000101",
    "1111010111110111",
    "1111000111111100",
    "1110111010010001",
    "1110110001001111",
    "1110101110110001",
    "1110110011111001",
    "1111000000001000",
    "1111010001111011",
    "1111100110111111",
    "1111111100111011",
    "1111101110101101",
    "1111011110001101",
    "1111010011011010",
    "1111001111011110",
    "1111010010111000",
    "1111011101001111",
    "1111101101101010",
    "1111111101010110",
    "1111100101110111",
    "1111001110011001",
    "1110111001101011",
    "1110101010001111",
    "1110100001111110",
    "1110100001101100",
    "1110101000111111",
    "1110110110010110",
    "1111000111011111",
    "1111011001101010",
    "1111101010000111",
    "1111110110010011",
    "1111111100001011",
    "1111111010100001",
    "1111110001001100",
    "1111100001010101",
    "1111001101001010",
    "1110110111100111",
    "1110100011100100",
    "1110010011011100",
    "1110001000011110",
    "1110000010110011",
    "1110000001011100",
    "1110000010111110",
    "1110000110000001",
    "1110001001101011",
    "1110001101101001",
    "1110010001110100",
    "1110010110010101",
    "1110011011010011",
    "1110100000111011",
    "1110100111011000",
    "1110101110111000",
    "1110110111101111",
    "1111000010100111",
    "1111010000010111",
    "1111100001101110",
    "1111110110111011",
    "1111110000110100",
    "1111010111100111",
    "1111000000001000",
    "1110101100111111",
    "1110011111110011",
    "1110011000101000",
    "1110010110001110",
    "1110010110100100",
    "1110010111101010",
    "1110011000100010",
    "1110011001101101",
    "1110011100111111",
    "1110100100101001",
    "1110110010000000",
    "1111000100101001",
    "1111011010001110",
    "1111101110111110",
    "1111111110110101",
    "1111111001010011",
    "1111111010111100",
    "1111111010011000",
    "1111101000110100",
    "1111010011011101",
    "1110111101110011",
    "1110101011001001",
    "1110011110000010",
    "1110011000001011",
    "1110011010010011",
    "1110100100011010",
    "1110110101110111",
    "1111001101000010",
    "1111100111001101",
    "1111111111001000",
    "1111101001110001",
    "1111011011100011",
    "1111010101101100",
    "1111010111101000",
    "1111011111010111",
    "1111101010010001",
    "1111110110001011",
    "1111111110001001",
    "1111110011000000",
    "1111100111111011",
    "1111011100010111",
    "1111010000010100",
    "1111000100101001",
    "1110111010111111",
    "1110110101010111",
    "1110110101101010",
    "1110111101000101",
    "1111001011100110",
    "1111011111111011",
    "1111110111101010",
    "1111110000000111",
    "1111011010011011",
    "1111001001101111",
    "1110111111101110",
    "1110111101001010",
    "1111000010000000",
    "1111001101101110",
    "1111011111101001",
    "1111110110110000",
    "1111101110011100",
    "1111010010001101",
    "1110110111001000",
    "1110011111110101",
    "1110001110010001",
    "1110000011100010",
    "1101111111011110",
    "1110000001001010",
    "1110000111000011",
    "1110001111100011",
    "1110011001011101",
    "1110100100000110",
    "1110101111100011",
    "1110111100001001",
    "1111001010010001",
    "1111011001101111",
    "1111101001100011",
    "1111110111111110",
    "1111111101000110",
    "1111110111011111",
    "1111111000000110",
    "1111111110101100",
    "1111110101111111",
    "1111101000000100",
    "1111011001111101",
    "1111001110001100",
    "1111000111001001",
    "1111000110111001",
    "1111001111001000",
    "1111100000011110",
    "1111111001111010",
    "1111100111011100",
    "1111001000000100",
    "1110101100110111",
    "1110011010000001",
    "1110010001110110",
    "1110010100001101",
    "1110011110110101",
    "1110101110001100",
    "1110111110101001",
    "1111001101100001",
    "1111011001011001",
    "1111100010111001",
    "1111101100101011",
    "1111111001111010",
    "1111110011011111",
    "1111011100000111",
    "1111000011000101",
    "1110101101000111",
    "1110011110111010",
    "1110011011100001",
    "1110100011000001",
    "1110110010100111",
    "1111000110000110",
    "1111011001010000",
    "1111101001001101",
    "1111110101000001",
    "1111111101001010",
    "1111111100111100",
    "1111110111110110",
    "1111110010110010",
    "1111101101101011",
    "1111101001000001",
    "1111100101011010",
    "1111100011010000",
    "1111100010100100",
    "1111100011011000",
    "1111100110001000",
    "1111101011101100",
    "1111110101000110",
    "1111111101000110",
    "1111101011011001",
    "1111010111001011",
    "1111000010101111",
    "1110110000100110",
    "1110100010111000",
    "1110011010101101",
    "1110010111111110",
    "1110011001100011",
    "1110011110001101",
    "1110100101010000",
    "1110101110111011",
    "1110111100000001",
    "1111001100110010",
    "1111100000011111",
    "1111110100111011",
    "1111111001001100",
    "1111101101000010",
    "1111101000011011",
    "1111101011010010",
    "1111110011100111",
    "1111111110100101",
    "1111110110011101",
    "1111101101001011",
    "1111100101111001",
    "1111100000000111",
    "1111011011001110",
    "1111010111010101",
    "1111010101010111",
    "1111010110111100",
    "1111011101101001",
    "1111101010000110",
    "1111111011100000",
    "1111110000011000",
    "1111011100110000",
    "1111001100110111",
    "1111000011010101",
    "1111000001101110",
    "1111001000011000",
    "1111010110100000",
    "1111101010011100",
    "1111111110001000",
    "1111100110000011",
    "1111001111111111",
    "1110111110000101",
    "1110110001100110",
    "1110101010110000",
    "1110101000111001",
    "1110101010111100",
    "1110101111111010",
    "1110110111000011",
    "1111000000000101",
    "1111001010101111",
    "1111010110011101",
    "1111100010001111",
    "1111101100110001",
    "1111110100110001",
    "1111111001011010",
    "1111111010101001",
    "1111111001000110",
    "1111110101111010",
    "1111110010001110",
    "1111101111000000",
    "1111101101000001",
    "1111101101000010",
    "1111101111111111",
    "1111110111000101",
    "1111111100101111",
    "1111101011100010",
    "1111010110101000",
    "1111000000100111",
    "1110101100101000",
    "1110011101011001",
    "1110010100011100",
    "1110010001101100",
    "1110010011110011",
    "1110011000111001",
    "1110011111011001",
    "1110100110100010",
    "1110101110011111",
    "1110110111111110",
    "1111000011110001",
    "1111010010011111",
    "1111100100010000",
    "1111111000101011",
    "1111110001001000",
    "1111011010110101",
    "1111000110100100",
    "1110110110101010",
    "1110101101000010",
    "1110101010101111",
    "1110101111011110",
    "1110111001101111",
    "1111000111001110",
    "1111010101111011",
    "1111100101000101",
    "1111110101010100",
    "1111111000000100",
    "1111100010100100",
    "1111001011001010",
    "1110110100110001",
    "1110100011010000",
    "1110011010000010",
    "1110011010110000",
    "1110100100011000",
    "1110110011101001",
    "1111000100010010",
    "1111010010010010",
    "1111011010111100",
    "1111011101010001",
    "1111011001101010",
    "1111010001010100",
    "1111000101111011",
    "1110111001000111",
    "1110101100101101",
    "1110100010010010",
    "1110011011011011",
    "1110011001011000",
    "1110011100110111",
    "1110100101111001",
    "1110110011101010",
    "1111000100101110",
    "1111010111001000",
    "1111101000111000",
    "1111111000001001",
    "1111111100100001",
    "1111110110001011",
    "1111110100111110",
    "1111111000010011",
    "1111111110110100",
    "1111111001010011",
    "1111110010001001",
    "1111101101011110",
    "1111101100011111",
    "1111101111101010",
    "1111110110101000",
    "1111111111100111",
    "1111110100101010",
    "1111101010000101",
    "1111100001010100",
    "1111011011001111",
    "1111011000001110",
    "1111010111111110",
    "1111011001111010",
    "1111011101011100",
    "1111100010000110",
    "1111100111101010",
    "1111101110000100",
    "1111110101011100",
    "1111111101110001",
    "1111111001010111",
    "1111110001000100",
    "1111101010110110",
    "1111101000011100",
    "1111101011011111",
    "1111110101000010",
    "1111111010111111",
    "1111100110001001",
    "1111001111001000",
    "1110111001001100",
    "1110100111011011",
    "1110011011111111",
    "1110010111100111",
    "1110011001110000",
    "1110100000111101",
    "1110101011011001",
    "1110110111100010",
    "1111000100010101",
    "1111010001001010",
    "1111011101110000",
    "1111101001101111",
    "1111110100100111",
    "1111111101101100",
    "1111111011100100",
    "1111110111100001",
    "1111110101111010",
    "1111110110000011",
    "1111110110111010",
    "1111110111100000",
    "1111110111001000",
    "1111110101100100",
    "1111110010110111",
    "1111101111001110",
    "1111101010110101",
    "1111100101110100",
    "1111100000010010",
    "1111011010010110",
    "1111010100001101",
    "1111001110001111",
    "1111001000111010",
    "1111000100101111",
    "1111000010011101",
    "1111000010110011",
    "1111000110100000",
    "1111001110000111",
    "1111011001110010",
    "1111101001000110",
    "1111111010111100",
    "1111110010010110",
    "1111100000110101",
    "1111010010010010",
    "1111000111111111",
    "1111000010100010",
    "1111000001101110",
    "1111000100110100",
    "1111001010110000",
    "1111010010100100",
    "1111011011011011",
    "1111100100110011",
    "1111101110100100",
    "1111111000111100",
    "1111111011011111",
    "1111101110001100",
    "1111011110110011",
    "1111001101110111",
    "1110111101000010",
    "1110101110110001",
    "1110100101100101",
    "1110100011010011",
    "1110101000100000",
    "1110110100101001",
    "1111000110010110",
    "1111011011110000",
    "1111110010100011",
    "1111110111101011",
    "1111100101011111",
    "1111011000110101",
    "1111010010111011",
    "1111010011111011",
    "1111011010101111",
    "1111100101101001",
    "1111110010110000",
    "1111111111011100",
    "1111110010000010",
    "1111100101101110",
    "1111011011001100",
    "1111010011010010",
    "1111001110110000",
    "1111001110000101",
    "1111010001000010",
    "1111010110100010",
    "1111011100101101",
    "1111100001010101",
    "1111100010100001",
    "1111011111010001",
    "1111010111110111",
    "1111001101101001",
    "1111000010011101",
    "1110111000000011",
    "1110101111101100",
    "1110101010000111",
    "1110100111011010",
    "1110100111010001",
    "1110101001011000",
    "1110101101010001",
    "1110110010011100",
    "1110111000010101",
    "1110111110001101",
    "1111000011010000",
    "1111000110110111",
    "1111001000110100",
    "1111001001100010",
    "1111001001111100",
    "1111001011010001",
    "1111001110101001",
    "1111010100110011",
    "1111011101111101",
    "1111101001111111",
    "1111111000110001",
    "1111110101111101",
    "1111100010111101",
    "1111001111100001",
    "1110111101100011",
    "1110101111001100",
    "1110100110000110",
    "1110100011001000",
    "1110100110000100",
    "1110101101111111",
    "1110111001100011",
    "1111000111111100",
    "1111011000110100",
    "1111101100010101",
    "1111111101110010",
    "1111100110110010",
    "1111010000110110",
    "1110111110110000",
    "1110110010111101",
    "1110101110110001",
    "1110110010000010",
    "1110111011001010",
    "1111000111110100",
    "1111010101110010",
    "1111100011101010",
    "1111110000111010",
    "1111111101010010",
    "1111110111100100",
    "1111101110101001",
    "1111101001001001",
    "1111101000001001",
    "1111101100000000",
    "1111110011110100",
    "1111111101101001",
    "1111111001000010",
    "1111110010101011",
    "1111110000110001",
    "1111110011110000",
    "1111111011001101",
    "1111111001110011",
    "1111101100100011",
    "1111011110010100",
    "1111010000011001",
    "1111000100000110",
    "1110111010100011",
    "1110110100100100",
    "1110110010100010",
    "1110110100010111",
    "1110111001101010",
    "1111000010001011",
    "1111001110000010",
    "1111011101100001",
    "1111110000101110",
    "1111111001001110",
    "1111100010010100",
    "1111001101001100",
    "1110111100100101",
    "1110110010010010",
    "1110101110110110",
    "1110110001011010",
    "1110111000001100",
    "1111000001011100",
    "1111001011111000",
    "1111010110111100",
    "1111100010100010",
    "1111101110100110",
    "1111111010110100",
    "1111111001010100",
    "1111101110100100",
    "1111100101100010",
    "1111011110101000",
    "1111011010000001",
    "1111010111101111",
    "1111010111101111",
    "1111011010000111",
    "1111011110111011",
    "1111100110001001",
    "1111101111001100",
    "1111111001000001",
    "1111111101101110",
    "1111110110011011",
    "1111110010000011",
    "1111110000111100",
    "1111110010101101",
    "1111110110011011",
    "1111111010111100",
    "1111111111100001",
    "1111111100000010",
    "1111110111011100",
    "1111110010001101",
    "1111101100000111",
    "1111100101101110",
    "1111100000011100",
    "1111011110010111",
    "1111100001100001",
    "1111101010110010",
    "1111111001011101",
    "1111110100110111",
    "1111100011101110",
    "1111010110100010",
    "1111001111111000",
    "1111010000110000",
    "1111011000101111",
    "1111100110100001",
    "1111111000110001",
    "1111110001010000",
    "1111011000010101",
    "1110111101011100",
    "1110100010100110",
    "1110001010010110",
    "1101110111010101",
    "1101101011010011",
    "1101100110100101",
    "1101101000000001",
    "1101101101001111",
    "1101110011110100",
    "1101111001111001",
    "1101111110101110",
    "1110000010011100",
    "1110000101101100",
    "1110001001010101",
    "1110001110001100",
    "1110010101001000",
    "1110011110111010",
    "1110101100001111",
    "1110111101000101",
    "1111010000101001",
    "1111100100111110",
    "1111110111011111",
    "1111111010011011",
    "1111110010110111",
    "1111110010100010",
    "1111111000110001",
    "1111111100000001",
    "1111101101110111",
    "1111011110110001",
    "1111010000100011",
    "1111000100101110",
    "1110111100100011",
    "1110111001000010",
    "1110111010110111",
    "1111000010001011",
    "1111001110011011",
    "1111011101111111",
    "1111101110101010",
    "1111111110000111",
    "1111110101100000",
    "1111101101000110",
    "1111101000011101",
    "1111100110101000",
    "1111100110100001",
    "1111100111011111",
    "1111101001101111",
    "1111101110010100",
    "1111110110110001",
    "1111111011101111",
    "1111101001001100",
    "1111010010111101",
    "1110111011111111",
    "1110100111111111",
    "1110011010100011",
    "1110010101111110",
    "1110011010110111",
    "1110101000001011",
    "1110111011111111",
    "1111010100000110",
    "1111101110100001",
    "1111110110101011",
    "1111011101110011",
    "1111001001001011",
    "1110111010111100",
    "1110110100100111",
    "1110110110100111",
    "1110111111111111",
    "1111001110110101",
    "1111100000111110",
    "1111110100100100",
    "1111110111110100",
    "1111100101010011",
    "1111010100110100",
    "1111000111010110",
    "1110111101110111",
    "1110111001001001",
    "1110111001100000",
    "1110111110100100",
    "1111000111100011",
    "1111010011101100",
    "1111100010010111",
    "1111110011011100",
    "1111111001001100",
    "1111100100000110",
    "1111001110101000",
    "1110111010111101",
    "1110101011101101",
    "1110100011000011",
    "1110100010000011",
    "1110101000010011",
    "1110110100001011",
    "1111000011010101",
    "1111010011010111",
    "1111100010011100",
    "1111101111011000",
    "1111111001110010",
    "1111111110011111",
    "1111111001011011",
    "1111110110111001",
    "1111110110101100",
    "1111111000011000",
    "1111111011010000",
    "1111111110011000",
    "1111111111000111",
    "1111111110000110",
    "1111111110111110",
    "1111111110000111",
    "1111111001010010",
    "1111110010100101",
    "1111101010000100",
    "1111011111110110",
    "1111010100010010",
    "1111001000000100",
    "1110111100010111",
    "1110110010011111",
    "1110101011101111",
    "1110101000111100",
    "1110101010010001",
    "1110101111001111",
    "1110110110110010",
    "1110111111110000",
    "1111001001001100",
    "1111010011100111",
    "1111100000110110",
    "1111110011000011",
    "1111110100111111",
    "1111011001000001",
    "1110111101001110",
    "1110100111001011",
    "1110011100011011",
    "1110100000010100",
    "1110110010010111",
    "1111001110001101",
    "1111101101001111",
    "1111110111011010",
    "1111100100101110",
    "1111011100101000",
    "1111011110011100",
    "1111100111011011",
    "1111110100011101",
    "1111111100101110",
    "1111101101001010",
    "1111011100110111",
    "1111001011101101",
    "1110111010100000",
    "1110101010101101",
    "1110011110000101",
    "1110010101111001",
    "1110010010010000",
    "1110010010011100",
    "1110010100110111",
    "1110010111111110",
    "1110011010100101",
    "1110011100011100",
    "1110011110001010",
    "1110100000110011",
    "1110100101100000",
    "1110101101001010",
    "1110111000001011",
    "1111000110010010",
    "1111010110010110",
    "1111100110100110",
    "1111110100101110",
    "1111111110101001",
    "1111111100110101",
    "1111111101110000",
    "1111111101001010",
    "1111110110010100",
    "1111110000001011",
    "1111101100100000",
    "1111101011110110",
    "1111101101011001",
    "1111101111101000",
    "1111110001000001",
    "1111110000011101",
    "1111101101101001",
    "1111101001000100",
    "1111100011110100",
    "1111011111010001",
    "1111011100100110",
    "1111011100101101",
    "1111011111111010",
    "1111100110001110",
    "1111101111001101",
    "1111111001110001",
    "1111111011101100",
    "1111110011001111",
    "1111101110110001",
    "1111101111111000",
    "1111110111011100",
    "1111111010100011",
    "1111100111011000",
    "1111010001001000",
    "1110111010011101",
    "1110100110000000",
    "1110010101111011",
    "1110001011011011",
    "1110000110110001",
    "1110000111010000",
    "1110001011100101",
    "1110010010010000",
    "1110011010000001",
    "1110100001111011",
    "1110101001011110",
    "1110110000011111",
    "1110110111000001",
    "1110111101001100",
    "1111000011000101",
    "1111001000011110",
    "1111001101000000",
    "1111010000000101",
    "1111010001001100",
    "1111001111111000",
    "1111001100000010",
    "1111000101110100",
    "1110111101110011",
    "1110110101000001",
    "1110101100110000",
    "1110100110100010",
    "1110100011110011",
    "1110100101100111",
    "1110101100011001",
    "1110110111100111",
    "1111000110000000",
    "1111010101101100",
    "1111100100101100",
    "1111110001010010",
    "1111111010010101",
    "1111111111011010",
    "1111111111001101",
    "1111111110111111",
    "1111111010110110",
    "1111110101000010",
    "1111101110001010",
    "1111100110101111",
    "1111011111010001",
    "1111011000001110",
    "1111010010001111",
    "1111001101110000",
    "1111001011010011",
    "1111001011001100",
    "1111001101101000",
    "1111010010101011",
    "1111011010011101",
    "1111100101001001",
    "1111110011001001",
    "1111111011000101",
    "1111100101101110",
    "1111001101110111",
    "1110110101101110",
    "1110100000000101",
    "1110001111101001",
    "1110000110001001",
    "1110000100000000",
    "1110001000010110",
    "1110010001100111",
    "1110011110101000",
    "1110101110111011",
    "1111000010010111",
    "1111011000010001",
    "1111101110110011",
    "1111111100111111",
    "1111101110101000",
    "1111101000111100",
    "1111101101000111",
    "1111111010000010",
    "1111110011010111",
    "1111011111010010",
    "1111001101101001",
    "1111000001011010",
    "1110111011111111",
    "1110111101010110",
    "1111000100011010",
    "1111001111011111",
    "1111011100100110",
    "1111101001101111",
    "1111110101001011",
    "1111111101100111",
    "1111111101101011",
    "1111111100110010",
    "1111111111000000",
    "1111111100110011",
    "1111111000000001",
    "1111110011110001",
    "1111110000110011",
    "1111101111010111",
    "1111101111010010",
    "1111110000001001",
    "1111110001011000",
    "1111110010010110",
    "1111110010100001",
    "1111110001011011",
    "1111101110100110",
    "1111101001100010",
    "1111100001110100",
    "1111010111010001",
    "1111001010100000",
    "1110111100101101",
    "1110101111100100",
    "1110100100101100",
    "1110011101000101",
    "1110011000111100",
    "1110010111100111",
    "1110010111111111",
    "1110011001000110",
    "1110011010100000",
    "1110011100110101",
    "1110100001101100",
    "1110101010111010",
    "1110111001011000",
    "1111001100011100",
    "1111100001100111",
    "1111110101000110",
    "1111111100110101",
    "1111110110110011",
    "1111111001001100",
    "1111111101100101",
    "1111110000010110",
    "1111100001111001",
    "1111010100010011",
    "1111001000100101",
    "1110111111001010",
    "1110111000010000",
    "1110110100011111",
    "1110110100101111",
    "1110111001111100",
    "1111000100011010",
    "1111010011101001",
    "1111100110000001",
    "1111111001011000",
    "1111110100011110",
    "1111100101001101",
    "1111011001100010",
    "1111010001011010",
    "1111001100011001",
    "1111001001101111",
    "1111001000110010",
    "1111001001000111",
    "1111001010100000",
    "1111001100111010",
    "1111010000011100",
    "1111010101001000",
    "1111011010110100",
    "1111100001000011",
    "1111100111001101",
    "1111101100011011",
    "1111110000000010",
    "1111110001101001",
    "1111110001001111",
    "1111101111010001",
    "1111101100100101",
    "1111101010010001",
    "1111101001101001",
    "1111101011110111",
    "1111110001110101",
    "1111111011111110",
    "1111110101111011",
    "1111100100110111",
    "1111010010010101",
    "1111000000010001",
    "1110110000100001",
    "1110100100101100",
    "1110011101101101",
    "1110011011110011",
    "1110011110101000",
    "1110100101011000",
    "1110101111000111",
    "1110111010110111",
    "1111000111111100",
    "1111010110000001",
    "1111100100111011",
    "1111110100100000",
    "1111111011101001",
    "1111101100101001",
    "1111011111110101",
    "1111010110101100",
    "1111010010011100",
    "1111010011100100",
    "1111011001110101",
    "1111100100100101",
    "1111110011000001",
    "1111111011011001",
    "1111100111100100",
    "1111010010101111",
    "1110111110110001",
    "1110101101111000",
    "1110100010000010",
    "1110011100100001",
    "1110011101100001",
    "1110100100010010",
    "1110101111010111",
    "1110111101010100",
    "1111001100111111",
    "1111011101001100",
    "1111101100101100",
    "1111111001110111",
    "1111111101000010",
    "1111111001100101",
    "1111111100010111",
    "1111111011010010",
    "1111101111011110",
    "1111100011001011",
    "1111011001100011",
    "1111010101000101",
    "1111010111000110",
    "1111011111011111",
    "1111101101000010",
    "1111111101101111",
    "1111110000100101",
    "1111100000000010",
    "1111010010001010",
    "1111000111110111",
    "1111000001011010",
    "1110111110100011",
    "1110111110011111",
    "1111000000001101",
    "1111000010100111",
    "1111000100110011",
    "1111000110001000",
    "1111000110100000",
    "1111000110001011",
    "1111000101101110",
    "1111000101110110",
    "1111000111010001",
    "1111001010100101",
    "1111010000000101",
    "1111011000000011",
    "1111100010101100",
    "1111110000010110",
    "1111111110110010",
    "1111101011001001",
    "1111010101110111",
    "1111000001000111",
    "1110101111010110",
    "1110100010110110",
    "1110011100110011",
    "1110011101001010",
    "1110100010110011",
    "1110101100010001",
    "1110111000101100",
    "1111001000010000",
    "1111011011110111",
    "1111110100000011",
    "1111110000000010",
    "1111010011010000",
    "1110111001100000",
    "1110100110011011",
    "1110011100011100",
    "1110011011110000",
    "1110100010101011",
    "1110101110101110",
    "1110111101111010",
    "1111001111011110",
    "1111100011100010",
    "1111111010001000",
    "1111101101110111",
    "1111010111001001",
    "1111000100111110",
    "1110111010010011",
    "1110111000011110",
    "1110111110110101",
    "1111001010110000",
    "1111011000111111",
    "1111100110101100",
    "1111110010001010",
    "1111111010111101",
    "1111111110101110",
    "1111111010101110",
    "1111111001001001",
    "1111111010010110",
    "1111111110101011",
    "1111111001111011",
    "1111110000010001",
    "1111100101100111",
    "1111011011100011",
    "1111010011011111",
    "1111001110101000",
    "1111001101111011",
    "1111010010011111",
    "1111011101100001",
    "1111101111111101",
    "1111110110100010",
    "1111011000001011",
    "1110111000011110",
    "1110011011110000",
    "1110000101101110",
    "1101111000100101",
    "1101110100100000",
    "1101110111110100",
    "1101111111111000",
    "1110001010010001",
    "1110010101011010",
    "1110100000101001",
    "1110101100000001",
    "1110111000001001",
    "1111000110010011",
    "1111010111111001",
    "1111101101100010",
    "1111111001011100",
    "1111011111010010",
    "1111000111001101",
    "1110110100101010",
    "1110101010011011",
    "1110101001100000",
    "1110110000110000",
    "1110111101010010",
    "1111001011110010",
    "1111011001010101",
    "1111100100010000",
    "1111101100000011",
    "1111110000111001",
    "1111110011000000",
    "1111110010010011",
    "1111101110011011",
    "1111100111010101",
    "1111011101101001",
    "1111010010111000",
    "1111001001010001",
    "1111000011000011",
    "1111000001101100",
    "1111000101010111",
    "1111001101000111",
    "1111010111001110",
    "1111100001110110",
    "1111101011110110",
    "1111110101100101",
    "1111111111011000",
    "1111110001011111",
    "1111100000010001",
    "1111001101001001",
    "1110111011000111",
    "1110101101111101",
    "1110101000101100",
    "1110101100100001",
    "1110111000010001",
    "1111001000111111",
    "1111011010111000",
    "1111101010100101",
    "1111110101110000",
    "1111111011011101",
    "1111111011110110",
    "1111110111111111",
    "1111110001010101",
    "1111101001011001",
    "1111100001100010",
    "1111011010110101",
    "1111010101110110",
    "1111010010110001",
    "1111010001010100",
    "1111010000110000",
    "1111010000001010",
    "1111001110110011",
    "1111001100010001",
    "1111001000101111",
    "1111000100100111",
    "1111000000011100",
    "1110111100111111",
    "1110111011000111",
    "1110111100000100",
    "1111000001001000",
    "1111001011100001",
    "1111011011110010",
    "1111110001001100",
    "1111110110000111",
    "1111011101001010",
    "1111000111001000",
    "1110110110011010",
    "1110101100000101",
    "1110100111101111",
    "1110100111101101",
    "1110101010000001",
    "1110101101000000",
    "1110101111111000",
    "1110110010111001",
    "1110110110101111",
    "1110111100001100",
    "1111000011100010",
    "1111001100011001",
    "1111010101101100",
    "1111011110000101",
    "1111100100010101",
    "1111100111100101",
    "1111100111101001",
    "1111100100111011",
    "1111100000010100",
    "1111011011000001",
    "1111010110010011",
    "1111010011011101",
    "1111010011100111",
    "1111010111101111",
    "1111100000101110",
    "1111101111011000",
    "1111111011110000",
    "1111100001000000",
    "1111000001111001",
    "1110100001100111",
    "1110000100010010",
    "1101101101110111",
    "1101100001001000",
    "1101011110110101",
    "1101100101100111",
    "1101110010111001",
    "1110000011111110",
    "1110010110111111",
    "1110101011011001",
    "1111000001010101",
    "1111011000110101",
    "1111110000111100",
    "1111111000011001",
    "1111100101101111",
    "1111011001010011",
    "1111010100000011",
    "1111010101100111",
    "1111011100011110",
    "1111100110111000",
    "1111110011100001",
    "1111111101111110",
    "1111101101101110",
    "1111011011111000",
    "1111001001100011",
    "1110111000110111",
    "1110101100010001",
    "1110100110000011",
    "1110100111011000",
    "1110101111111000",
    "1110111101110010",
    "1111001110010010",
    "1111011110011110",
    "1111101011110010",
    "1111110100100010",
    "1111110111111110",
    "1111110110001011",
    "1111101111111001",
    "1111100110011000",
    "1111011011000100",
    "1111001111100100",
    "1111000101010011",
    "1110111101010110",
    "1110111000001011",
    "1110110101110100",
    "1110110101111011",
    "1110111000000001",
    "1110111011101111",
    "1111000000111011",
    "1111000111101101",
    "1111010000010100",
    "1111011010110100",
    "1111100111010101",
    "1111110101110000",
    "1111111010001100",
    "1111101001011100",
    "1111011001011000",
    "1111001100000010",
    "1111000011011111",
    "1111000001110000",
    "1111001000001100",
    "1111010111011101",
    "1111101110110111",
    "1111110011110100",
    "1111010100010010",
    "1110110110110010",
    "1110011111011001",
    "1110010000110110",
    "1110001100000010",
    "1110001111110110",
    "1110011001101010",
    "1110100110011101",
    "1110110011110001",
    "1111000000001010",
    "1111001011010001",
    "1111010101001000",
    "1111011101111000",
    "1111100101010011",
    "1111101010111101",
    "1111101110010111",
    "1111101111100010",
    "1111101111000110",
    "1111101110011000",
    "1111101110111011",
    "1111110001111010",
    "1111110111110100",
    "1111111111101011",
    "1111110101100111",
    "1111101011001100",
    "1111100001100100",
    "1111011001100111",
    "1111010011110011",
    "1111010000001010",
    "1111001110100100",
    "1111001110101001",
    "1111010000000010",
    "1111010010001011",
    "1111010100101001",
    "1111010110110100",
    "1111011000001011",
    "1111011000010001",
    "1111010110111011",
    "1111010100010000",
    "1111010000101100",
    "1111001100111000",
    "1111001001011011",
    "1111000110111001",
    "1111000101110010",
    "1111000110101000",
    "1111001001111111",
    "1111010000011001",
    "1111011001111010",
    "1111100110000011",
    "1111110011011011",
    "1111111111110010",
    "1111110101100100",
    "1111101111010111",
    "1111101101110011",
    "1111110000100100",
    "1111110110100011",
    "1111111110010101",
    "1111111001011000",
    "1111110001101000",
    "1111101010100110",
    "1111100011110011",
    "1111011100001100",
    "1111010011000000",
    "1111001000010101",
    "1110111101011100",
    "1110110100100100",
    "1110110000001111",
    "1110110010011001",
    "1110111011100001",
    "1111001010101000",
    "1111011101010001",
    "1111110000100001",
    "1111111110001110",
    "1111110000101110",
    "1111100111100101",
    "1111100010011100",
    "1111100000011111",
    "1111100000110001",
    "1111100010101100",
    "1111100101110111",
    "1111101010010000",
    "1111101111101111",
    "1111110110000100",
    "1111111100110101",
    "1111111100011011",
    "1111110110001111",
    "1111110000111110",
    "1111101100110111",
    "1111101010000000",
    "1111101000001011",
    "1111100110110111",
    "1111100101001110",
    "1111100010010101",
    "1111011101001111",
    "1111010101011000",
    "1111001010101010",
    "1110111101100001",
    "1110101110111010",
    "1110011111111011",
    "1110010001101011",
    "1110000100111001",
    "1101111010001001",
    "1101110001101100",
    "1101101011110101",
    "1101101000111111",
    "1101101001110000",
    "1101101110100110",
    "1101110111100101",
    "1110000100010010",
    "1110010011101001",
    "1110100100010111",
    "1110110101000110",
    "1111000100111011",
    "1111010011001010",
    "1111011111011111",
    "1111101001110101",
    "1111110001111001",
    "1111110111011000",
    "1111111010000010",
    "1111111001111000",
    "1111110111010110",
    "1111110011001100",
    "1111101110010010",
    "1111101001001100",
    "1111100100001000",
    "1111011110110110",
    "1111011000111111",
    "1111010010100001",
    "1111001011111111",
    "1111000110101000",
    "1111000100000011",
    "1111000101100010",
    "1111001011101101",
    "1111010110000000",
    "1111100010101111",
    "1111101111100101",
    "1111111010000001",
    "1111111111111110",
    "1111111111110010",
    "1111111010001110",
    "1111101110101110",
    "1111011111010010",
    "1111001110010001",
    "1110111110010100",
    "1110110001111110",
    "1110101011001100",
    "1110101010110101",
    "1110110000110001",
    "1110111100000001",
    "1111001011000100",
    "1111011100011011",
    "1111101110110101",
    "1111111110110100",
    "1111101101100111",
    "1111011110100100",
    "1111010010100111",
    "1111001010010001",
    "1111000101100111",
    "1111000100000000",
    "1111000100011000",
    "1111000101100101",
    "1111000110101100",
    "1111000111010101",
    "1111000111101100",
    "1111001000011010",
    "1111001010000100",
    "1111001101001010",
    "1111010001111001",
    "1111011000010001",
    "1111100000010100",
    "1111101010000010",
    "1111110101011101",
    "1111111101100000",
    "1111101111101011",
    "1111100010010000",
    "1111010110110100",
    "1111001110110001",
    "1111001010110101",
    "1111001010111010",
    "1111001110000010",
    "1111010010111101",
    "1111011000100101",
    "1111011110101011",
    "1111100101101110",
    "1111101110110010",
    "1111111010110011",
    "1111110110001010",
    "1111100101010000",
    "1111010100101111",
    "1111000111100000",
    "1111000000001000",
    "1111000000010010",
    "1111001000011000",
    "1111010111101010",
    "1111101100010111",
    "1111111100000110",
    "1111100100110001",
    "1111010000011111",
    "1111000001100111",
    "1110111001100000",
    "1110111000001001",
    "1110111100010011",
    "1111000011111011",
    "1111001100111101",
    "1111010101101110",
    "1111011101011011",
    "1111100100000000",
    "1111101001111000",
    "1111101111100000",
    "1111110101001001",
    "1111111010101110",
    "1111111111111011",
    "1111111011100011",
    "1111110111111100",
    "1111110101000110",
    "1111110010101110",
    "1111110000100001",
    "1111101110010010",
    "1111101011111011",
    "1111101001010011",
    "1111100110001001",
    "1111100010000011",
    "1111011100100101",
    "1111010101010111",
    "1111001100010110",
    "1111000010000000",
    "1110110111001000",
    "1110101100111000",
    "1110100100100101",
    "1110011111010001",
    "1110011101100001",
    "1110011111100001",
    "1110100100110100",
    "1110101100101101",
    "1110110110010110",
    "1111000000111011",
    "1111001011110010",
    "1111010110010101",
    "1111100000010010",
    "1111101001011110",
    "1111110001111011",
    "1111111001101101",
    "1111111111000111",
    "1111111000110101",
    "1111110011101110",
    "1111110000000111",
    "1111101110010001",
    "1111101110010001",
    "1111110000000010",
    "1111110011010110",
    "1111110111111000",
    "1111111101010011",
    "1111111100110000",
    "1111110110110100",
    "1111110001011100",
    "1111101101010011",
    "1111101011000111",
    "1111101011010101",
    "1111101110000001",
    "1111110010101011",
    "1111111000011000",
    "1111111101111001",
    "1111111101111000",
    "1111111011111011",
    "1111111100100100",
    "1111111111110101",
    "1111111010011100",
    "1111110010011011",
    "1111101000001000",
    "1111011011101000",
    "1111001101010111",
    "1110111110011100",
    "1110110000100111",
    "1110100101110111",
    "1110011111110000",
    "1110011110111000",
    "1110100010011101",
    "1110101000110010",
    "1110101111101000",
    "1110110101000000",
    "1110110111110100",
    "1110110111111110",
    "1110110110000110",
    "1110110011001011",
    "1110110000001100",
    "1110101101110011",
    "1110101100011100",
    "1110101100001001",
    "1110101100110010",
    "1110101110000111",
    "1110101111101011",
    "1110110001000000",
    "1110110001011111",
    "1110110000100100",
    "1110101101111111",
    "1110101001101111",
    "1110100100010011",
    "1110011110100100",
    "1110011001100011",
    "1110010110011010",
    "1110010110000110",
    "1110011001010011",
    "1110100000011010",
    "1110101011100011",
    "1110111010101010",
    "1111001101100001",
    "1111100011100111",
    "1111111011111011",
    "1111101011010101",
    "1111010100101110",
    "1111000010100010",
    "1110110110100010",
    "1110110001001111",
    "1110110001101110",
    "1110110110010010",
    "1110111100111111",
    "1111000100110001",
    "1111001101111000",
    "1111011001101000",
    "1111101001100110",
    "1111111110001111",
    "1111101001110011",
    "1111010001110011",
    "1110111101101001",
    "1110110000100110",
    "1110101100000100",
    "1110101111001100",
    "1110110111011010",
    "1111000001100001",
    "1111001010110101",
    "1111010001110110",
    "1111010110000110",
    "1111010111110010",
    "1111010111001000",
    "1111010100010000",
    "1111001111010001",
    "1111001000011010",
    "1111000000011001",
    "1110111000011000",
    "1110110001110110",
    "1110101110001100",
    "1110101110011100",
    "1110110011001000",
    "1110111100010011",
    "1111001001110000",
    "1111011011010100",
    "1111110000101110",
    "1111110110110100",
    "1111011100111010",
    "1111000011101111",
    "1110101101101001",
    "1110011100011011",
    "1110010000110110",
    "1110001010100010",
    "1110001000011000",
    "1110001000111110",
    "1110001011010110",
    "1110001111010110",
    "1110010101010011",
    "1110011101110011",
    "1110101000111111",
    "1110110110001110",
    "1111000100001010",
    "1111010000110001",
    "1111011010001110",
    "1111011111010010",
    "1111011111101001",
    "1111011011111000",
    "1111010101000101",
    "1111001100011100",
    "1111000011001011",
    "1110111010001100",
    "1110110010010100",
    "1110101100000101",
    "1110101000000100",
    "1110100110100101",
    "1110100111111010",
    "1110101100001110",
    "1110110011100111",
    "1110111110001111",
    "1111001011111101",
    "1111011100001111",
    "1111101101111111",
    "1111111111011001",
    "1111110001100001",
    "1111100110101000",
    "1111100000111001",
    "1111100000011010",
    "1111100100011010",
    "1111101011101010",
    "1111110101001100",
    "1111111111000110",
    "1111110000111010",
    "1111100000000011",
    "1111001101011100",
    "1110111011001111",
    "1110101100001010",
    "1110100010110100",
    "1110100000101100",
    "1110100101110100",
    "1110110000111001",
    "1111000000010001",
    "1111010010011100",
    "1111100110010110",
    "1111111010111010",
    "1111110001011011",
    "1111100001000000",
    "1111010110011000",
    "1111010011101110",
    "1111011010000110",
    "1111101000101111",
    "1111111101001011",
    "1111101100000110",
    "1111010110111110",
    "1111000110100010",
    "1110111100101101",
    "1110111010000111",
    "1110111110011100",
    "1111001000101000",
    "1111010111010011",
    "1111101000101010",
    "1111111010110100",
    "1111110011111010",
    "1111100100111001",
    "1111011000101000",
    "1111001110111000",
    "1111000110110001",
    "1110111111011010",
    "1110111000010001",
    "1110110001011100",
    "1110101011100011",
    "1110100111011000",
    "1110100101100100",
    "1110100110001101",
    "1110101001000001",
    "1110101101010100",
    "1110110010011010",
    "1110110111110101",
    "1110111101100001",
    "1111000011110100",
    "1111001011001110",
    "1111010100000011",
    "1111011110010010",
    "1111101001100000",
    "1111110101000000",
    "1111111111110110",
    "1111110101110100",
    "1111101101011010",
    "1111100111001100",
    "1111100011101110",
    "1111100011011111",
    "1111100110100111",
    "1111101100101010",
    "1111110100011111",
    "1111111100011111",
    "1111111100111110",
    "1111111001010000",
    "1111111000111001",
    "1111111011110101",
    "1111111110010011",
    "1111110101111111",
    "1111101011010110",
    "1111011110100011",
    "1111010000001100",
    "1111000001011111",
    "1110110100011000",
    "1110101011000100",
    "1110100111011000",
    "1110101010010011",
    "1110110011101010",
    "1111000010001011",
    "1111010011111110",
    "1111100110110111",
    "1111111000101110",
    "1111111000001111",
    "1111101101100000",
    "1111101000000010",
    "1111101000010100",
    "1111101110010101",
    "1111111001100001",
    "1111110111000111",
    "1111100101001101",
    "1111010010011010",
    "1111000000011110",
    "1110110000110000",
    "1110100100000011",
    "1110011010101101",
    "1110010100101111",
    "1110010010001000",
    "1110010011000110",
    "1110011000000001",
    "1110100001011100",
    "1110101111100001",
    "1111000001111001",
    "1111010111010001",
    "1111101101101100",
    "1111111101010001",
    "1111101011111101",
    "1111011111111011",
    "1111011001110111",
    "1111011001010110",
    "1111011101001111",
    "1111100100000001",
    "1111101100001110",
    "1111110100100011",
    "1111111100001000",
    "1111111101100001",
    "1111111000101001",
    "1111110101001101",
    "1111110011001100",
    "1111110010101101",
    "1111110011111010",
    "1111110110111100",
    "1111111011101110",
    "1111111110000100",
    "1111110111001011",
    "1111110000100100",
    "1111101011010011",
    "1111101000011001",
    "1111101000100101",
    "1111101100010111",
    "1111110100000100",
    "1111111111111101",
    "1111101111100111",
    "1111011011000111",
    "1111000011111000",
    "1110101100001111",
    "1110010111011000",
    "1110001000010000",
    "1110000000111110",
    "1110000010001010",
    "1110001010110010",
    "1110011000111110",
    "1110101010111000",
    "1110111111101000",
    "1111010110111111",
    "1111110000110010",
    "1111110011111000",
    "1111011001010001",
    "1111000010100010",
    "1110110011001000",
    "1110101101101011",
    "1110110010111011",
    "1111000001100001",
    "1111010110001011",
    "1111101100110000",
    "1111111110101110",
    "1111101111011000",
    "1111100110110101",
    "1111100101100010",
    "1111101011000001",
    "1111110110000100",
    "1111111011000011",
    "1111101010100101",
    "1111011010110010",
    "1111001101101110",
    "1111000100110001",
    "1111000000011001",
    "1111000000000011",
    "1111000010011111",
    "1111000110010101",
    "1111001010100110",
    "1111001110111011",
    "1111010011010101",
    "1111011000000110",
    "1111011101010110",
    "1111100010111011",
    "1111101000011010",
    "1111101101010001",
    "1111110001000101",
    "1111110011101111",
    "1111110101011000",
    "1111110110010001",
    "1111110110101011",
    "1111110110101110",
    "1111110110011100",
    "1111110101111011",
    "1111110101011010",
    "1111110101001110",
    "1111110101101100",
    "1111110110111000",
    "1111111000100011",
    "1111111010000011",
    "1111111010100100",
    "1111111001011101",
    "1111110110100000",
    "1111110010001000",
    "1111101101010001",
    "1111101001000101",
    "1111100110110010",
    "1111100111011000",
    "1111101011100011",
    "1111110011111000",
    "1111111111001100",
    "1111101101111000",
    "1111011001010001",
    "1111000011011111",
    "1110101111011100",
    "1110011111111111",
    "1110010111001011",
    "1110010101101001",
    "1110011010011000",
    "1110100011011000",
    "1110101110011011",
    "1110111001111001",
    "1111000101001110",
    "1111010000101011",
    "1111011100110011",
    "1111101001110101",
    "1111110111010000",
    "1111111100000111",
    "1111110001111100",
    "1111101011011101",
    "1111101001010001",
    "1111101011000000",
    "1111101111100101",
    "1111110101100101",
    "1111111011100111",
    "1111111111011100",
    "1111111100100000",
    "1111111100000111",
    "1111111110101100",
    "1111111011100001",
    "1111110010101100",
    "1111100111010100",
    "1111011010011110",
    "1111001101110000",
    "1111000010111001",
    "1110111011100011",
    "1110111000111010",
    "1110111011101000",
    "1111000011100111",
    "1111010000001010",
    "1111100000000011",
    "1111110001101101",
    "1111111100101011",
    "1111101100111011",
    "1111100000010101",
    "1111010111100111",
    "1111010010101111",
    "1111010001001000",
    "1111010001111000",
    "1111010100001010",
    "1111010111011111",
    "1111011011101010",
    "1111100000110101",
    "1111100111010000",
    "1111101111000100",
    "1111111000001000",
    "1111111101111001",
    "1111110011101100",
    "1111101001111000",
    "1111100001010000",
    "1111011010101010",
    "1111010110111110",
    "1111010111000100",
    "1111011011101010",
    "1111100100110110",
    "1111110001111100",
    "1111111110011010",
    "1111101110011101",
    "1111100000011110",
    "1111010110011011",
    "1111010001101011",
    "1111010010011111",
    "1111011000010011",
    "1111100001111011",
    "1111101110000100",
    "1111111011101010",
    "1111110110000111",
    "1111101000000111",
    "1111011011010100",
    "1111010001000111",
    "1111001010111111",
    "1111001010001011",
    "1111001110110110",
    "1111011000000011",
    "1111100011011111",
    "1111101110010000",
    "1111110101011110",
    "1111110111000101",
    "1111110010000101",
    "1111100110100111",
    "1111010101110010",
    "1111000001100110",
    "1110101100010001",
    "1110011000010000",
    "1110000111100010",
    "1101111011011110",
    "1101110100101100",
    "1101110010111110",
    "1101110101101100",
    "1101111011111010",
    "1110000100111001",
    "1110010000001100",
    "1110011101010111",
    "1110101100000100",
    "1110111011101011",
    "1111001011001110",
    "1111011001100111",
    "1111100101110010",
    "1111101111001011",
    "1111110101101101",
    "1111111001111010",
    "1111111100110000",
    "1111111111010011",
    "1111111101100001",
    "1111111001010000",
    "1111110011110000",
    "1111101101001110",
    "1111100110001000",
    "1111011111000010",
    "1111011000101000",
    "1111010011011101",
    "1111001111111111",
    "1111001110011100",
    "1111001110111101",
    "1111010001110100",
    "1111011000010001",
    "1111100100010010",
    "1111110111100101",
    "1111101101101111",
    "1111001110010001",
    "1110101110101001",
    "1110010100010111",
    "1110000011111011",
    "1101111111010100",
    "1110000101001011",
    "1110010001101110",
    "1110100000010101",
    "1110101101101101",
    "1110111001000001",
    "1111000011100001",
    "1111001111010110",
    "1111011101111010",
    "1111101110110100",
    "1111111111111000",
    "1111110010001100",
    "1111101010011100",
    "1111101010001111",
    "1111110000110111",
    "1111111011110111",
    "1111110111110000",
    "1111101100100110",
    "1111100100001010",
    "1111011110111111",
    "1111011101000100",
    "1111011101111101",
    "1111100001001111",
    "1111100110011101",
    "1111101101001001",
    "1111110100101110",
    "1111111100010010",
    "1111111101001101",
    "1111111000111001",
    "1111110111100111",
    "1111111001110101",
    "1111111111101110",
    "1111110110111111",
    "1111101011001001",
    "1111011101110111",
    "1111010000101011",
    "1111000101010011",
    "1110111101010110",
    "1110111001111001",
    "1110111011001111",
    "1111000000111011",
    "1111001001110111",
    "1111010100110100",
    "1111100000110000",
    "1111101100111100",
    "1111111000111111",
    "1111111011010100",
    "1111110000000111",
    "1111100101011101",
    "1111011011011110",
    "1111010010011100",
    "1111001010100110",
    "1111000100011100",
    "1111000000010101",
    "1110111110111101",
    "1111000001000010",
    "1111000111000011",
    "1111010001000101",
    "1111011110011001",
    "1111101101011110",
    "1111111100010011",
    "1111110111001100",
    "1111101110110001",
    "1111101011001110",
    "1111101100011010",
    "1111110001011001",
    "1111111000111001",
    "1111111110000111",
    "1111110100010011",
    "1111101001111100",
    "1111011111011110",
    "1111010101101100",
    "1111001110000010",
    "1111001010001111",
    "1111001100000010",
    "1111010100010111",
    "1111100010101100",
    "1111110100111001",
    "1111111000011100",
    "1111101001001011",
    "1111100000010010",
    "1111011111010100",
    "1111100110000011",
    "1111110010100011",
    "1111111101110110",
    "1111101101111000",
    "1111011111011001",
    "1111010011010111",
    "1111001001111101",
    "1111000011001011",
    "1110111110111011",
    "1110111101010110",
    "1110111110101011",
    "1111000010111110",
    "1111001001111001",
    "1111010010101100",
    "1111011100010110",
    "1111100101110100",
    "1111101110011101",
    "1111110110001000",
    "1111111101010000",
    "1111111011100010",
    "1111110011110010",
    "1111101011010100",
    "1111100010011101",
    "1111011001111010",
    "1111010010100111",
    "1111001101011011",
    "1111001010111101",
    "1111001011010100",
    "1111001110000111",
    "1111010010100010",
    "1111010111101010",
    "1111011100100110",
    "1111100001010100",
    "1111100110111100",
    "1111101111111100",
    "1111111110110100",
    "1111101010111000",
    "1111001110000000",
    "1110101101110011",
    "1110001110111010",
    "1101110110001001",
    "1101100110101010",
    "1101100000111011",
    "1101100011000001",
    "1101101001100101",
    "1101110001010101",
    "1101111000100101",
    "1101111111010001",
    "1110000110011010",
    "1110001110110110",
    "1110011000010101",
    "1110100000111011",
    "1110100101111100",
    "1110100100110111",
    "1110011100111000",
    "1110001111100001",
    "1110000000001100",
    "1101110011000011",
    "1101101011011000",
    "1101101010100101",
    "1101110000011111",
    "1101111100001100",
    "1110001101010010",
    "1110100011101110",
    "1110111111001100",
    "1111011110001101",
    "1111111101101110",
    "1111100110010011",
    "1111010001110011",
    "1111000110111111",
    "1111000101011111",
    "1111001010100000",
    "1111010010010111",
    "1111011001111101",
    "1111100000001101",
    "1111100101111011",
    "1111101100111010",
    "1111110110110100",
    "1111111100000000",
    "1111101100111111",
    "1111011110101110",
    "1111010100001010",
    "1111001111011110",
    "1111010001100111",
    "1111011010000110",
    "1111100111010010",
    "1111110111001000",
    "1111111000101001",
    "1111101010010000",
    "1111011111010110",
    "1111011000110101",
    "1111010110110111",
    "1111011000101010",
    "1111011100111010",
    "1111100010000011",
    "1111100110111000",
    "1111101010101101",
    "1111101101100101",
    "1111110000000000",
    "1111110010100011",
    "1111110101100011",
    "1111111000111011",
    "1111111100010001",
    "1111111111000110",
    "1111111110111011",
    "1111111101110101",
    "1111111101010110",
    "1111111101000100",
    "1111111100110111",
    "1111111100111110",
    "1111111101110011",
    "1111111111101010",
    "1111111101100001",
    "1111111010011100",
    "1111111000001011",
    "1111111000000111",
    "1111111011100110",
    "1111111100010111",
    "1111101111101100",
    "1111011111011111",
    "1111001110000010",
    "1110111110001010",
    "1110110010101011",
    "1110101101011110",
    "1110101111001101",
    "1110110111000011",
    "1111000011010000",
    "1111010001111110",
    "1111100001110110",
    "1111110010011011",
    "1111111100011100",
    "1111101011010010",
    "1111011011001110",
    "1111001110001101",
    "1111000110010110",
    "1111000101001101",
    "1111001010111111",
    "1111010110010011",
    "1111100100011000",
    "1111110010001010",
    "1111111100111111",
    "1111111100011010",
    "1111111010000100",
    "1111111010110011",
    "1111111100111001",
    "1111111110101000",
    "1111111110101110",
    "1111111100101000",
    "1111111000011001",
    "1111110010101111",
    "1111101100101011",
    "1111100111010111",
    "1111100011110100",
    "1111100010111000",
    "1111100100111001",
    "1111101001110011",
    "1111110001001101",
    "1111111010011010",
    "1111111011011101",
    "1111110001011101",
    "1111101000011110",
    "1111100001010101",
    "1111011100101011",
    "1111011010111100",
    "1111011100100001",
    "1111100001101011",
    "1111101010001011",
    "1111110101010110",
    "1111111110000010",
    "1111110001101001",
    "1111100111000111",
    "1111011111101100",
    "1111011011111000",
    "1111011011011101",
    "1111011101100110",
    "1111100001011010",
    "1111100110010010",
    "1111101100000011",
    "1111110010111100",
    "1111111011001011",
    "1111111011001001",
    "1111110000101001",
    "1111100110011111",
    "1111011110011111",
    "1111011010110010",
    "1111011101000111",
    "1111100110001110",
    "1111110101100000",
    "1111110111000111",
    "1111100010110100",
    "1111010000111101",
    "1111000100010011",
    "1110111110100110",
    "1111000000001010",
    "1111001000011000",
    "1111010110010010",
    "1111101001000010",
    "1111111111111001",
    "1111100101010000",
    "1111001000011010",
    "1110101011110010",
    "1110010010011100",
    "1101111111011100",
    "1101110100110011",
    "1101110010111011",
    "1101111000101010",
    "1110000011110100",
    "1110010001111011",
    "1110100001000000",
    "1110101111101000",
    "1110111100111100",
    "1111001000001110",
    "1111010000110011",
    "1111010101111110",
    "1111010111010000",
    "1111010100100010",
    "1111001110011001",
    "1111000101110111",
    "1110111100010111",
    "1110110011010101",
    "1110101100000101",
    "1110100111101101",
    "1110100111000100",
    "1110101010110010",
    "1110110011001101",
    "1111000000000111",
    "1111010000011111",
    "1111100010101111",
    "1111110100110001",
    "1111111011011001",
    "1111101111001110",
    "1111100111010001",
    "1111100011011000",
    "1111100010110110",
    "1111100100110001",
    "1111101000011011",
    "1111101101010010",
    "1111110011000000",
    "1111111001010101",
    "1111111111111110",
    "1111111001001000",
    "1111110010000100",
    "1111101010100001",
    "1111100010000000",
    "1111011000001100",
    "1111001101011100",
    "1111000010110100",
    "1110111010000111",
    "1110110101001001",
    "1110110101010010",
    "1110111010111111",
    "1111000101111001",
    "1111010100110111",
    "1111100110011000",
    "1111111000100100",
    "1111110110101000",
    "1111101001010101",
    "1111100001001100",
    "1111011111010010",
    "1111100100000000",
    "1111101110111100",
    "1111111111010011",
    "1111101100000111",
    "1111010101001101",
    "1110111110010001",
    "1110101010000100",
    "1110011011000010",
    "1110010010111001",
    "1110010001110110",
    "1110010110110010",
    "1110011111011110",
    "1110101001010000",
    "1110110001110001",
    "1110110111100111",
    "1110111010010001",
    "1110111010000110",
    "1110110111101111",
    "1110110100000001",
    "1110101111100001",
    "1110101010101000",
    "1110100101110001",
    "1110100001011100",
    "1110011110010111",
    "1110011101001010",
    "1110011110001101",
    "1110100001100001",
    "1110100110110110",
    "1110101101110010",
    "1110110101111100",
    "1110111111000100",
    "1111001000111110",
    "1111010011011111",
    "1111011110101001",
    "1111101010011101",
    "1111110111000010",
    "1111111011100001",
    "1111101101011001",
    "1111011110111000",
    "1111010000100001",
    "1111000011000001",
    "1110110111001001",
    "1110101101011100",
    "1110100110001000",
    "1110100001000011",
    "1110011101110010",
    "1110011011110010",
    "1110011010101000",
    "1110011010001100",
    "1110011010110101",
    "1110011101001001",
    "1110100001111110",
    "1110101010010100",
    "1110110110111110",
    "1111001000000100",
    "1111011100110000",
    "1111110011000001",
    "1111111000000111",
    "1111100111110111",
    "1111011110101011",
    "1111011101011100",
    "1111100011010010",
    "1111101101110011",
    "1111111001111010",
    "1111111011001001",
    "1111110011010001",
    "1111101111000010",
    "1111101110000010",
    "1111101111010101",
    "1111110001111010",
    "1111110101000110",
    "1111111000011010",
    "1111111011011101",
    "1111111101110100",
    "1111111110110110",
    "1111111101111001",
    "1111111010011111",
    "1111110100011100",
    "1111101100000000",
    "1111100001111001",
    "1111010111000110",
    "1111001100101110",
    "1111000011110100",
    "1110111101000101",
    "1110111000110010",
    "1110110110101111",
    "1110110110010110",
    "1110110110111110",
    "1110111000000110",
    "1110111001101000",
    "1110111011101010",
    "1110111110011110",
    "1111000010001011",
    "1111000110011111",
    "1111001010110010",
    "1111001110000111",
    "1111001111100110",
    "1111001110101011",
    "1111001011100000",
    "1111000110110010",
    "1111000001111110",
    "1110111110110101",
    "1110111111000000",
    "1111000011101110",
    "1111001101001001",
    "1111011010001111",
    "1111101001000010",
    "1111110111000111",
    "1111111101011110",
    "1111110101110110",
    "1111110001110010",
    "1111110000001001",
    "1111101111011101",
    "1111101110100001",
    "1111101100110011",
    "1111101010010110",
    "1111100111100000",
    "1111100100100010",
    "1111100001011111",
    "1111011110000111",
    "1111011010001111",
    "1111010101111001",
    "1111010001011111",
    "1111001101101101",
    "1111001011010100",
    "1111001011000110",
    "1111001101100011",
    "1111010011000011",
    "1111011011101011",
    "1111100111001111",
    "1111110101000111",
    "1111111011110100",
    "1111101101010110",
    "1111100001011010",
    "1111011001110111",
    "1111010111111010",
    "1111011011100110",
    "1111100011101100",
    "1111101101111000",
    "1111110111010100",
    "1111111101001110",
    "1111111101100110",
    "1111110111100001",
    "1111101011011100",
    "1111011011000010",
    "1111001000111001",
    "1110110111101111",
    "1110101001111100",
    "1110100001001000",
    "1110011101111010",
    "1110100000010001",
    "1110100111100111",
    "1110110011010111",
    "1111000010110100",
    "1111010101010011",
    "1111101001100110",
    "1111111110000011",
    "1111101111011000",
    "1111100000101110",
    "1111010111010000",
    "1111010011001011",
    "1111010011100111",
    "1111010110110001",
    "1111011010101101",
    "1111011101110011",
    "1111011111001111",
    "1111011111000111",
    "1111011110001100",
    "1111011101100110",
    "1111011110010110",
    "1111100001001101",
    "1111100110100011",
    "1111101110011000",
    "1111111000011110",
    "1111111011010110",
    "1111101101010100",
    "1111011101100110",
    "1111001100101101",
    "1110111011110000",
    "1110101100000111",
    "1110011111001100",
    "1110010110000011",
    "1110010001000000",
    "1110001111101011",
    "1110010001000101",
    "1110010100001011",
    "1110011000011010",
    "1110011101111011",
    "1110100101101010",
    "1110110000101110",
    "1110111111101110",
    "1111010010001010",
    "1111100110001110",
    "1111111000111111",
    "1111111000101100",
    "1111110001011100",
    "1111110010011100",
    "1111111011010100",
    "1111110101100111",
    "1111100011001000",
    "1111010000001010",
    "1110111111100100",
    "1110110011100010",
    "1110101101001111",
    "1110101100110010",
    "1110110001010000",
    "1110111001000111",
    "1111000010101001",
    "1111001100010011",
    "1111010101000001",
    "1111011100011001",
    "1111100010100001",
    "1111100111110010",
    "1111101100101001",
    "1111110001011000",
    "1111110110000010",
    "1111111010011101",
    "1111111110011110",
    "1111111101111110",
    "1111111010111010",
    "1111111000000111",
    "1111110101011100",
    "1111110010110011",
    "1111110000000101",
    "1111101101001010",
    "1111101001110110",
    "1111100101111011",
    "1111100001001111",
    "1111011011111010",
    "1111010110010010",
    "1111010000111001",
    "1111001100010111",
    "1111001001001011",
    "1111000111100111",
    "1111000111101010",
    "1111001000111100",
    "1111001010111111",
    "1111001101100100",
    "1111010000110000",
    "1111010100110111",
    "1111011010100010",
    "1111100010010000",
    "1111101100010111",
    "1111111000101000",
    "1111111001100110",
    "1111101011100100",
    "1111011110101101",
    "1111010100011010",
    "1111001101110010",
    "1111001011011000",
    "1111001101010110",
    "1111010011100110",
    "1111011110000010",
    "1111101100010011",
    "1111111101100001",
    "1111101111110011",
    "1111011101110101",
    "1111001110101110",
    "1111000100001110",
    "1110111111001111",
    "1110111111011110",
    "1111000011111100",
    "1111001011010011",
    "1111010100001010",
    "1111011101010111",
    "1111100101101111",
    "1111101011111000",
    "1111101110001010",
    "1111101011000000",
    "1111100001011010",
    "1111010001101110",
    "1110111101111010",
    "1110101001001100",
    "1110010111001110",
    "1110001011001001",
    "1110000110101111",
    "1110001010000111",
    "1110010100001000",
    "1110100011000001",
    "1110110101000000",
    "1111001000011010",
    "1111011011111000",
    "1111101110000001",
    "1111111101011010",
    "1111110111010101",
    "1111110001010000",
    "1111110000101001",
    "1111110100110101",
    "1111111100001101",
    "1111111011011011",
    "1111110100010110",
    "1111110000010001",
    "1111110000000001",
    "1111110011011011",
    "1111111001011011",
    "1111111111100000",
    "1111111001000010",
    "1111110100011100",
    "1111110010100100",
    "1111110011101111",
    "1111110111101100",
    "1111111101111100",
    "1111111010001111",
    "1111110001110000",
    "1111101001100010",
    "1111100010101001",
    "1111011110000101",
    "1111011100110101",
    "1111011111011110",
    "1111100110010101",
    "1111110001001111",
    "1111111111011111",
    "1111110000001000",
    "1111011111010111",
    "1111010000000000",
    "1111000011100010",
    "1110111010111000",
    "1110110110000100",
    "1110110100011101",
    "1110110101000011",
    "1110110110111110",
    "1110111001111111",
    "1110111110100001",
    "1111000101011010",
    "1111001111010111",
    "1111011100010100",
    "1111101011001001",
    "1111111001100111",
    "1111111011000011",
    "1111110101011011",
    "1111110110110010",
    "1111111110101001",
    "1111110101000100",
    "1111100111100000",
    "1111011011110000",
    "1111010100001011",
    "1111010001110001",
    "1111010100011000",
    "1111011011000100",
    "1111100100110001",
    "1111110000101111",
    "1111111110011101",
    "1111110010100010",
    "1111100011001011",
    "1111010100110111",
    "1111001001001110",
    "1111000001110100",
    "1110111111101100",
    "1111000010111101",
    "1111001011000100",
    "1111010110111111",
    "1111100101011111",
    "1111110101010010",
    "1111111010101111",
    "1111101011111010",
    "1111011111010001",
    "1111010101101100",
    "1111001111110000",
    "1111001101101101",
    "1111001111011111",
    "1111010100110100",
    "1111011101010100",
    "1111101000011010",
    "1111110101011100",
    "1111111100010110",
    "1111101110000001",
    "1111100000101001",
    "1111010101010000",
    "1111001100101110",
    "1111000111101100",
    "1111000110010010",
    "1111001000010110",
    "1111001101100001",
    "1111010101010000",
    "1111011110111010",
    "1111101001101110",
    "1111110100110110",
    "1111111111010011",
    "1111110111111001",
    "1111110001101111",
    "1111101110110010",
    "1111101111010011",
    "1111110011001100",
    "1111111010001100",
    "1111111100000010",
    "1111101111111000",
    "1111100001111101",
    "1111010011010111",
    "1111000101101111",
    "1110111011000010",
    "1110110101000110",
    "1110110101001000",
    "1110111011100110",
    "1111001000001000",
    "1111011001101101",
    "1111101110110111",
    "1111111010100111",
    "1111100101011111",
    "1111010100100111",
    "1111001010100011",
    "1111001000111010",
    "1111010000001100",
    "1111011111111011",
    "1111110111000101",
    "1111101011111011",
    "1111001011100110",
    "1110101011001001",
    "1110001110010010",
    "1101111000100010",
    "1101101100001111",
    "1101101010001011",
    "1101110001010101",
    "1101111111011110",
    "1110010001101100",
    "1110100101011111",
    "1110111000111010",
    "1111001010110000",
    "1111011010001111",
    "1111100110110111",
    "1111110000001010",
    "1111110101111000",
    "1111111000000100",
    "1111110111010111",
    "1111110101000011",
    "1111110010101100",
    "1111110001110001",
    "1111110011000110",
    "1111110110101010",
    "1111111011110000",
    "1111111110101010",
    "1111111001110010",
    "1111110110100000",
    "1111110101100010",
    "1111110111001110",
    "1111111011100000",
    "1111111110000001",
    "1111110110001111",
    "1111101110000001",
    "1111100110010101",
    "1111011111111011",
    "1111011011100000",
    "1111011001011001",
    "1111011001110010",
    "1111011100011100",
    "1111100000111110",
    "1111100110101111",
    "1111101101000011",
    "1111110011000111",
    "1111111000001000",
    "1111111011010011",
    "1111111011110011",
    "1111111001000100",
    "1111110010111011",
    "1111101001111001",
    "1111011111001010",
    "1111010100011100",
    "1111001011100000",
    "1111000101111110",
    "1111000100110001",
    "1111001000001000",
    "1111001111101100",
    "1111011010111101",
    "1111101001101000",
    "1111111011110000",
    "1111101110101011",
    "1111010110101010",
    "1110111110001010",
    "1110101000000011",
    "1110010111001011",
    "1110001101100110",
    "1110001100000100",
    "1110010001111000",
    "1110011101011001",
    "1110101100111000",
    "1110111111000100",
    "1111010011001000",
    "1111101000011010",
    "1111111101110111",
    "1111101110000100",
    "1111011101100001",
    "1111010010010100",
    "1111001101100100",
    "1111001111010001",
    "1111010110001011",
    "1111100000011110",
    "1111101100000001",
    "1111110111001010",
    "1111111111001100",
    "1111110111111001",
    "1111110011011011",
    "1111110010010000",
    "1111110100100111",
    "1111111010001110",
    "1111111101101100",
    "1111110100010110",
    "1111101011000010",
    "1111100010111011",
    "1111011100110010",
    "1111011000111111",
    "1111010111110001",
    "1111011001001001",
    "1111011101010010",
    "1111100100001011",
    "1111101101100100",
    "1111111000100111",
    "1111111011110100",
    "1111110001010010",
    "1111101001000110",
    "1111100100001110",
    "1111100011000101",
    "1111100101011011",
    "1111101010101111",
    "1111110010011010",
    "1111111011111001",
    "1111111001010011",
    "1111101101110001",
    "1111100010010100",
    "1111010111111001",
    "1111001111101001",
    "1111001010011101",
    "1111001000110100",
    "1111001010101010",
    "1111001111011010",
    "1111010110001101",
    "1111011110000010",
    "1111100110001110",
    "1111101110111110",
    "1111111001100111",
    "1111110111110111",
    "1111100100000011",
    "1111001011000010",
    "1110101111001000",
    "1110010100011000",
    "1101111111001100",
    "1101110010111011",
    "1101110000101001",
    "1101110110110110",
    "1110000010010000",
    "1110001111000010",
    "1110011001111101",
    "1110100000111101",
    "1110100010111101",
    "1110011111110011",
    "1110010111111111",
    "1110001100101010",
    "1101111111101001",
    "1101110011010101",
    "1101101010000001",
    "1101100101011111",
    "1101100110011010",
    "1101101100001110",
    "1101110101001000",
    "1101111111011111",
    "1110001011101000",
    "1110011011111000",
    "1110110010101001",
    "1111010000011001",
    "1111110010011010",
    "1111101100100110",
    "1111010010100111",
    "1111000100001101",
    "1111000010011100",
    "1111001010010100",
    "1111010110100111",
    "1111100001111011",
    "1111101000111101",
    "1111101011001100",
    "1111101010001111",
    "1111101000011111",
    "1111101000001000",
    "1111101001111111",
    "1111101101101100",
    "1111110010011001",
    "1111110111011111",
    "1111111101001101",
    "1111111011010010",
    "1111110000110110",
    "1111100011000101",
    "1111010010101110",
    "1111000001100110",
    "1110110001101100",
    "1110100100101110",
    "1110011011110010",
    "1110010111010001",
    "1110010110110111",
    "1110011001111010",
    "1110011111101001",
    "1110100111100111",
    "1110110001110011",
    "1110111110010001",
    "1111001100111101",
    "1111011101001110",
    "1111101101110000",
    "1111111100100110",
    "1111111000100001",
    "1111110011110000",
    "1111110110010011",
    "1111111111110001",
    "1111101111111000",
    "1111011100101011",
    "1111001001100000",
    "1110111001101010",
    "1110101111011111",
    "1110101011111101",
    "1110101110110000",
    "1110110110110110",
    "1111000011000110",
    "1111010010101100",
    "1111100100110100",
    "1111111000011110",
    "1111110011110100",
    "1111100001111110",
    "1111010011101110",
    "1111001010011110",
    "1111000110101111",
    "1111000111110101",
    "1111001100010100",
    "1111010010100001",
    "1111011000111100",
    "1111011110101001",
    "1111100011001010",
    "1111100110001001",
    "1111100111011010",
    "1111100110101000",
    "1111100011100001",
    "1111011110000101",
    "1111010110101111",
    "1111001110010100",
    "1111000101111011",
    "1110111110110011",
    "1110111010000110",
    "1110111000110111",
    "1110111011111100",
    "1111000011101110",
    "1111001111111011",
    "1111011111100011",
    "1111110001000110",
    "1111111101000010",
    "1111101100010000",
    "1111011101001110",
    "1111001111111011",
    "1111000011111011",
    "1110111000110111",
    "1110101110110011",
    "1110100110010000",
    "1110100000001100",
    "1110011101011100",
    "1110011110010111",
    "1110100010011111",
    "1110101000101111",
    "1110101111110001",
    "1110110110011010",
    "1110111100001001",
    "1111000001001100",
    "1111000110010010",
    "1111001100001110",
    "1111010011011101",
    "1111011011110111",
    "1111100100100010",
    "1111101100011001",
    "1111110010011000",
    "1111110101111010",
    "1111110111001011",
    "1111110110111110",
    "1111110110100100",
    "1111110111010000",
    "1111111010001001",
    "1111111111111011",
    "1111110111000110",
    "1111101011000110",
    "1111011100010100",
    "1111001011100000",
    "1110111001111001",
    "1110101001100010",
    "1110011100110101",
    "1110010110010010",
    "1110010111101010",
    "1110100001110001",
    "1110110011110011",
    "1111001011001111",
    "1111100100011100",
    "1111111011010111",
    "1111110011010001",
    "1111101001011111",
    "1111100111100111",
    "1111101100011100",
    "1111110101111101",
    "1111111101111100",
    "1111110001000110",
    "1111100100101001",
    "1111011001011000",
    "1111001111110101",
    "1111001000100101",
    "1111000100000000",
    "1111000010000110",
    "1111000010011100",
    "1111000011111100",
    "1111000101010000",
    "1111000100110110",
    "1111000001011010",
    "1110111010010100",
    "1110101111110101",
    "1110100011000011",
    "1110010101110001",
    "1110001001101011",
    "1110000000010100",
    "1101111010101010",
    "1101111000111111",
    "1101111011010001",
    "1110000001010010",
    "1110001010111010",
    "1110011000010001",
    "1110101001010110",
    "1110111101101001",
    "1111010100000000",
    "1111101010010101",
    "1111111110000100",
    "1111110011000111",
    "1111101010110010",
    "1111101001000100",
    "1111101100111011",
    "1111110100100111",
    "1111111110011101",
    "1111110110100011",
    "1111101010101011",
    "1111011101101011",
    "1111001111100110",
    "1111000001010100",
    "1110110100100111",
    "1110101011101010",
    "1110101000011000",
    "1110101011100110",
    "1110110100101110",
    "1111000001100110",
    "1111001111010111",
    "1111011011001010",
    "1111100010110011",
    "1111100100111110",
    "1111100001101011",
    "1111011001101101",
    "1111001110101101",
    "1111000010101011",
    "1110110111100101",
    "1110101111001100",
    "1110101010100101",
    "1110101010000111",
    "1110101101011110",
    "1110110011111000",
    "1110111100011001",
    "1111000110010010",
    "1111010000111101",
    "1111011100000001",
    "1111100111000101",
    "1111110001100101",
    "1111111010101100",
    "1111111110011110",
    "1111111010110011",
    "1111111010101111",
    "1111111110010011",
    "1111111010111011",
    "1111110001110101",
    "1111100111010101",
    "1111011100011001",
    "1111010001111001",
    "1111001000101000",
    "1111000001001010",
    "1110111011111111",
    "1110111001010011",
    "1110111001000111",
    "1110111011000100",
    "1110111110011100",
    "1111000010011100",
    "1111000110001101",
    "1111001001000110",
    "1111001010111101",
    "1111001011111111",
    "1111001100101101",
    "1111001101100110",
    "1111001111001000",
    "1111010001011100",
    "1111010100100000",
    "1111011000010000",
    "1111011100100110",
    "1111100001100111",
    "1111100111011001",
    "1111101110000001",
    "1111110101010100",
    "1111111100111101",
    "1111111011100010",
    "1111110100101000",
    "1111101110011000",
    "1111101000100011",
    "1111100010011111",
    "1111011011001111",
    "1111010001110011",
    "1111000101100111",
    "1110110111000011",
    "1110100111011111",
    "1110011000111010",
    "1110001101100011",
    "1110000110111110",
    "1110000101101111",
    "1110001001011000",
    "1110010000100110",
    "1110011010001011",
    "1110100101100000",
    "1110110010110110",
    "1111000010100111",
    "1111010100101110",
    "1111101000000010",
    "1111111010010110",
    "1111110111000010",
    "1111101110100000",
    "1111101101000101",
    "1111110010000100",
    "1111111011001010",
    "1111111010101000",
    "1111110010001110",
    "1111101101010111",
    "1111101100011101",
    "1111101110101110",
    "1111110010101010",
    "1111110110011110",
    "1111111000100111",
    "1111110111111100",
    "1111110011110011",
    "1111101100001001",
    "1111100001100100",
    "1111010101010111",
    "1111001001011001",
    "1110111111111000",
    "1110111010101111",
    "1110111011010001",
    "1111000001111101",
    "1111001110010001",
    "1111011110110101",
    "1111110001011011",
    "1111111100100001",
    "1111101101101000",
    "1111100011111110",
    "1111100000101110",
    "1111100100000101",
    "1111101101010010",
    "1111111011000000",
    "1111110100010000",
    "1111100001111000",
    "1111001110111010",
    "1110111100100000",
    "1110101011110101",
    "1110011110001010",
    "1110010100101110",
    "1110010000011100",
    "1110010001110100",
    "1110011000111010",
    "1110100101011011",
    "1110110110100101",
    "1111001011000010",
    "1111100000110110",
    "1111110101011011",
    "1111111001101011",
    "1111101110100101",
    "1111101010001010",
    "1111101100001100",
    "1111110011010011",
    "1111111101110010",
    "1111110101110100",
    "1111101000100100",
    "1111011010111010",
    "1111001101010111",
    "1111000000111011",
    "1110110111010001",
    "1110110010100100",
    "1110110100110011",
    "1110111110111010",
    "1111010000010100",
    "1111100110110000",
    "1111111110110110",
    "1111101010110111",
    "1111011001001100",
    "1111001101100001",
    "1111000111110010",
    "1111000111000011",
    "1111001010000001",
    "1111001111011111",
    "1111010110110010",
    "1111011111100011",
    "1111101001101001",
    "1111110100110110",
    "1111111111001111",
    "1111110011011110",
    "1111101000110100",
    "1111100000001101",
    "1111011010011001",
    "1111010111111100",
    "1111011000111111",
    "1111011101010111",
    "1111100100100100",
    "1111101101101110",
    "1111110111101010",
    "1111111110110000",
    "1111110110110001",
    "1111110001000110",
    "1111101110001100",
    "1111101101111111",
    "1111110000000111",
    "1111110011111111",
    "1111111000111110",
    "1111111110011010",
    "1111111100010000",
    "1111110111100001",
    "1111110011011111",
    "1111110000000100",
    "1111101100111100",
    "1111101001110001",
    "1111100110011011",
    "1111100011000101",
    "1111100000010100",
    "1111011110110011",
    "1111011111001100",
    "1111100001111000",
    "1111100110101111",
    "1111101101001011",
    "1111110100001010",
    "1111111010010110",
    "1111111110010111",
    "1111111111000110",
    "1111111011110010",
    "1111110100000110",
    "1111100111111000",
    "1111010111011011",
    "1111000011101001",
    "1110101110010110",
    "1110011010000001",
    "1110001001010001",
    "1101111110010110",
    "1101111010011000",
    "1101111101010100",
    "1110000110000011",
    "1110010011001111",
    "1110100100000000",
    "1110111000000011",
    "1111001111000010",
    "1111101000000000",
    "1111111110111111",
    "1111101000110001",
    "1111011000010000",
    "1111001111100001",
    "1111001111000111",
    "1111010101100101",
    "1111100000001101",
    "1111101011110001",
    "1111110101011010",
    "1111111011010100",
    "1111111100110110",
    "1111111010010010",
    "1111110100100010",
    "1111101100101110",
    "1111100100000101",
    "1111011011101011",
    "1111010100100000",
    "1111001111000111",
    "1111001011101010",
    "1111001001110111",
    "1111001001000110",
    "1111001000101000",
    "1111001000000100",
    "1111000111010011",
    "1111000110101100",
    "1111000110110001",
    "1111001000000100",
    "1111001010111100",
    "1111001111011010",
    "1111010101011000",
    "1111011100100110",
    "1111100101000110",
    "1111101111000100",
    "1111111010110010",
    "1111110111101001",
    "1111101000111011",
    "1111011010011001",
    "1111001101111000",
    "1111000101000101",
    "1111000000111101",
    "1111000001100110",
    "1111000101111100",
    "1111001100100011",
    "1111010011111000",
    "1111011010111100",
    "1111100001010101",
    "1111100111000101",
    "1111101100010101",
    "1111110000111111",
    "1111110100101110",
    "1111110110111100",
    "1111110110111101",
    "1111110100001000",
    "1111101110001110",
    "1111100101100000",
    "1111011010110101",
    "1111001111011111",
    "1111000100111110",
    "1110111100111000",
    "1110111000101100",
    "1110111001100000",
    "1111000000001111",
    "1111001101010110",
    "1111100000010111",
    "1111110111101110",
    "1111101111001110",
    "1111010111110111",
    "1111000101001000",
    "1110111000110101",
    "1110110011000101",
    "1110110010010100",
    "1110110100000110",
    "1110110110001000",
    "1110110110110111",
    "1110110110000001",
    "1110110100010010",
    "1110110010110100",
    "1110110010100010",
    "1110110011111100",
    "1110110110110110",
    "1110111010101010",
    "1110111110101001",
    "1111000010000010",
    "1111000100010011",
    "1111000101001000",
    "1111000100011000",
    "1111000010010010",
    "1110111111010010",
    "1110111100010011",
    "1110111010010100",
    "1110111010011110",
    "1110111101100100",
    "1111000100001000",
    "1111001110010100",
    "1111011100000010",
    "1111101100110011",
    "1111111111101011",
    "1111101100101000",
    "1111011001110010",
    "1111001001010001",
    "1110111100001100",
    "1110110011000000",
    "1110101101100011",
    "1110101011001110",
    "1110101011001110",
    "1110101100101110",
    "1110101111000111",
    "1110110001110011",
    "1110110100011100",
    "1110110110111001",
    "1110111001100010",
    "1110111101101000",
    "1111000100111110",
    "1111010001001111",
    "1111100010110100",
    "1111111000010101",
    "1111110001001110",
    "1111011101111101",
    "1111010001100110",
    "1111001110011100",
    "1111010100100101",
    "1111100010000101",
    "1111110011101011",
    "1111111010001001",
    "1111101010101010",
    "1111100000001111",
    "1111011100010011",
    "1111011111011010",
    "1111101001011000",
    "1111111001000011",
    "1111110011101001",
    "1111011111101100",
    "1111001110010001",
    "1111000010010000",
    "1110111101101001",
    "1111000001001000",
    "1111001100001001",
    "1111011101000100",
    "1111110001010111",
    "1111111001110101",
    "1111100111100011",
    "1111011010000001",
    "1111010010011010",
    "1111010000101011",
    "1111010011100010",
    "1111011001010000",
    "1111100000000010",
    "1111100110110111",
    "1111101101100001",
    "1111110100010110",
    "1111111011110100",
    "1111111011111010",
    "1111110011011010",
    "1111101011101000",
    "1111100101110111",
    "1111100011001000",
    "1111100100000000",
    "1111101000010010",
    "1111101111001101",
    "1111110111101011",
    "1111111111010000",
    "1111110110011100",
    "1111101110010100",
    "1111100111001101",
    "1111100001001111",
    "1111011100100001",
    "1111011001000110",
    "1111010110111100",
    "1111010110000011",
    "1111010110011000",
    "1111010111110001",
    "1111011001111101",
    "1111011100101011",
    "1111011111100100",
    "1111100010100111",
    "1111100101110110",
    "1111101001101001",
    "1111101110100000",
    "1111110100111100",
    "1111111101010111",
    "1111111000000000",
    "1111101011011001",
    "1111011101011011",
    "1111001111010100",
    "1111000010101111",
    "1110111001100010",
    "1110110101001101",
    "1110110110100101",
    "1110111101100100",
    "1111001001000100",
    "1111010111001001",
    "1111100101011111",
    "1111110001110100",
    "1111111010100011",
    "1111111111000001",
    "1111111111011110",
    "1111111100111110",
    "1111111001000010",
    "1111110101001011",
    "1111110010100101",
    "1111110001110101",
    "1111110010110100",
    "1111110100110101",
    "1111110110111100",
    "1111111000001010",
    "1111110111101101",
    "1111110101001111",
    "1111110000110111",
    "1111101011000000",
    "1111100100001110",
    "1111011100111111",
    "1111010101100111",
    "1111001110010001",
    "1111000110111110",
    "1110111111101110",
    "1110111000100010",
    "1110110001011010",
    "1110101010011011",
    "1110100011100100",
    "1110011100110010",
    "1110010101111100",
    "1110001111001000",
    "1110001000100101",
    "1110000010110011",
    "1101111110100110",
    "1101111100110101",
    "1101111110010100",
    "1110000011011100",
    "1110001100001001",
    "1110010111110010",
    "1110100101010101",
    "1110110011100110",
    "1111000001011110",
    "1111001110001100",
    "1111011001011000",
    "1111100010111011",
    "1111101010111101",
    "1111110001100101",
    "1111110110110011",
    "1111111010011100",
    "1111111100010000",
    "1111111100000010",
    "1111111001110011",
    "1111110101110100",
    "1111110000100001",
    "1111101010100011",
    "1111100100100101",
    "1111011111001100",
    "1111011010110111",
    "1111011000000100",
    "1111010111001001",
    "1111011000100111",
    "1111011100101101",
    "1111100011100111",
    "1111101101001100",
    "1111111000101000",
    "1111111011011110",
    "1111110001001110",
    "1111101010110100",
    "1111101010010011",
    "1111110001000011",
    "1111111111001001",
    "1111101100111101",
    "1111010110011011",
    "1111000001001000",
    "1110110000110101",
    "1110101000001001",
    "1110101000001011",
    "1110110000011010",
    "1110111111010100",
    "1111010011010010",
    "1111101011001001",
    "1111111010001000",
    "1111011110000111",
    "1111000011000001",
    "1110101011101011",
    "1110011010101011",
    "1110010001110000",
    "1110010001001000",
    "1110010111100111",
    "1110100011001000",
    "1110110001101011",
    "1111000001110011",
    "1111010010110011",
    "1111100100010011",
    "1111110101101011",
    "1111111010000111",
    "1111101100100000",
    "1111100010101111",
    "1111011101011011",
    "1111011100010011",
    "1111011110010001",
    "1111100001110000",
    "1111100101011000",
    "1111101000010100",
    "1111101010011000",
    "1111101011110101",
    "1111101101000101",
    "1111101110010110",
    "1111101111101011",
    "1111110001000100",
    "1111110010100011",
    "1111110100010111",
    "1111110111000101",
    "1111111011011010",
    "1111111101110101",
    "1111110100001101",
    "1111100111101000",
    "1111011000100011",
    "1111001000001011",
    "1110111000001011",
    "1110101010100000",
    "1110100001001101",
    "1110011101111000",
    "1110100001011111",
    "1110101011111000",
    "1110111011100101",
    "1111001110000010",
    "1111100000001100",
    "1111101111010111",
    "1111111001111100",
    "1111111111101110",
    "1111111110001111",
    "1111111110011000",
    "1111111111001001",
    "1111111111110000",
    "1111111111101110",
    "1111111110110110",
    "1111111101000100",
    "1111111010001110",
    "1111110110110001",
    "1111110011011111",
    "1111110001010000",
    "1111110000100101",
    "1111110001100001",
    "1111110011110000",
    "1111110110110100",
    "1111111010001110",
    "1111111101101000",
    "1111111111000111",
    "1111111100010001",
    "1111111010000110",
    "1111111001000011",
    "1111111001101100",
    "1111111100101000",
    "1111111101100100",
    "1111110100100110",
    "1111101000010110",
    "1111011001001100",
    "1111001000000110",
    "1110110110100000",
    "1110100110010000",
    "1110011001000111",
    "1110010000100011",
    "1110001101001110",
    "1110001111000010",
    "1110010101001000",
    "1110011110001100",
    "1110101000101111",
    "1110110011100010",
    "1110111101101011",
    "1111000110110001",
    "1111001110101011",
    "1111010101100100",
    "1111011011101010",
    "1111100001000011",
    "1111100101101010",
    "1111101001001110",
    "1111101011011100",
    "1111101011111001",
    "1111101010011001",
    "1111100111000001",
    "1111100010001000",
    "1111011100100000",
    "1111010110111110",
    "1111010010011101",
    "1111001111101001",
    "1111001110110011",
    "1111001111110011",
    "1111010010000011",
    "1111010100110100",
    "1111010111001110",
    "1111011000011011",
    "1111010111100101",
    "1111010011111011",
    "1111001100101000",
    "1111000001001111",
    "1110110010000110",
    "1110100000100110",
    "1110001111000010",
    "1110000000001100",
    "1101110110011010",
    "1101110011001101",
    "1101110110101100",
    "1101111111100011",
    "1110001011110111",
    "1110011001111010",
    "1110101001001001",
    "1110111010000010",
    "1111001101010110",
    "1111100011000101",
    "1111111001110101",
    "1111110001000010",
    "1111100000111000",
    "1111011000011011",
    "1111011000110010",
    "1111100000111000",
    "1111101101110011",
    "1111111011110110",
    "1111111000011000",
    "1111110001010000",
    "1111101111101011",
    "1111110011001110",
    "1111111010011011",
    "1111111100100100",
    "1111110011110001",
    "1111101100101001",
    "1111101000000111",
    "1111100110100101",
    "1111100111111100",
    "1111101011100110",
    "1111110000100100",
    "1111110101100100",
    "1111111001010111",
    "1111111011000100",
    "1111111010000111",
    "1111110110011110",
    "1111110000100100",
    "1111101001001010",
    "1111100001010010",
    "1111011010000001",
    "1111010100010010",
    "1111010000110000",
    "1111001111110000",
    "1111010001011010",
    "1111010101100100",
    "1111011100001010",
    "1111100101001110",
    "1111110000100111",
    "1111111101110010",
    "1111110100010001",
    "1111100111001000",
    "1111011100001010",
    "1111010100010111",
    "1111010000000010",
    "1111001110110001",
    "1111001111110000",
    "1111010001111110",
    "1111010100111100",
    "1111011000100010",
    "1111011100111100",
    "1111100010000011",
    "1111100111010010",
    "1111101011010110",
    "1111101100101001",
    "1111101001110100",
    "1111100010010111",
    "1111010110111001",
    "1111001001000110",
    "1110111011010011",
    "1110101111110110",
    "1110101000101000",
    "1110100110101000",
    "1110101010001111",
    "1110110011010111",
    "1111000001100110",
    "1111010100011010",
    "1111101011001001",
    "1111111011001001",
    "1111100000000010",
    "1111000101100000",
    "1110101101111011",
    "1110011011011011",
    "1110001111010100",
    "1110001001111010",
    "1110001010011110",
    "1110001111110011",
    "1110011000100010",
    "1110100011101001",
    "1110110000100110",
    "1110111110111111",
    "1111001110010010",
    "1111011101100001",
    "1111101011010101",
    "1111110110010000",
    "1111111101001000",
    "1111111111011100",
    "1111111101011001",
    "1111110111110100",
    "1111110000000101",
    "1111100111110000",
    "1111100000011110",
    "1111011011101011",
    "1111011010100110",
    "1111011101111011",
    "1111100101101010",
    "1111110000111110",
    "1111111110011100",
    "1111110011101010",
    "1111100111000110",
    "1111011101000111",
    "1111010110010110",
    "1111010011000000",
    "1111010010110001",
    "1111010101001110",
    "1111011010000111",
    "1111100001100001",
    "1111101100000010",
    "1111111010100001",
    "1111110010001010",
    "1111011001111101",
    "1110111110000111",
    "1110100001010111",
    "1110000111011101",
    "1101110011111110",
    "1101101001001110",
    "1101100111101010",
    "1101101101111000",
    "1101111001001001",
    "1110000110011101",
    "1110010011100111",
    "1110100000010001",
    "1110101101101001",
    "1110111101100110",
    "1111010001000101",
    "1111100111001110",
    "1111111101011000",
    "1111110000010001",
    "1111100101011010",
    "1111100100000110",
    "1111101100001101",
    "1111111011100100",
    "1111110001000100",
    "1111011101000100",
    "1111001011000110",
    "1110111101001010",
    "1110110100100101",
    "1110110001111101",
    "1110110101001011",
    "1110111101100011",
    "1111001001011101",
    "1111010110101100",
    "1111100010101111",
    "1111101011011101",
    "1111101111010110",
    "1111101110001110",
    "1111101001000010",
    "1111100001011010",
    "1111011000111111",
    "1111010001010000",
    "1111001011001100",
    "1111000111011101",
    "1111000110100000",
    "1111001000011000",
    "1111001100110101",
    "1111010011001010",
    "1111011010001110",
    "1111100000110001",
    "1111100101101111",
    "1111101000011011",
    "1111101000100011",
    "1111100110010011",
    "1111100010010000",
    "1111011101001100",
    "1111011000000100",
    "1111010011111011",
    "1111010001011010",
    "1111010000111001",
    "1111010010011001",
    "1111010101011010",
    "1111011001010001",
    "1111011101000100",
    "1111100000000000",
    "1111100001100010",
    "1111100001011100",
    "1111011111101100",
    "1111011100100001",
    "1111011000000100",
    "1111010010011101",
    "1111001011101111",
    "1111000011111100",
    "1110111011001100",
    "1110110001110011",
    "1110101000010001",
    "1110011111100001",
    "1110011000100000",
    "1110010100001110",
    "1110010011010111",
    "1110010110010011",
    "1110011101010001",
    "1110101000011110",
    "1110111000001011",
    "1111001100010001",
    "1111100011111100",
    "1111111101100100",
    "1111101001011000",
    "1111010011111001",
    "1111000100011111",
    "1110111100101000",
    "1110111100001100",
    "1111000001100001",
    "1111001001111001",
    "1111010010010010",
    "1111010111111111",
    "1111011001010000",
    "1111010101100100",
    "1111001101100100",
    "1111000010110110",
    "1110110111010001",
    "1110101100101000",
    "1110100100001010",
    "1110011110100011",
    "1110011011111010",
    "1110011011110010",
    "1110011101010111",
    "1110011111110110",
    "1110100010100010",
    "1110100101010011",
    "1110101000110111",
    "1110101111010001",
    "1110111011001010",
    "1111001110100100",
    "1111101001100000",
    "1111110110011110",
    "1111010110000011",
    "1110111010011110",
    "1110101000001100",
    "1110100001010000",
    "1110100100110001",
    "1110101111110101",
    "1110111110110110",
    "1111001111000000",
    "1111011110111000",
    "1111101110010001",
    "1111111101101100",
    "1111110010010111",
    "1111100010010000",
    "1111010011000110",
    "1111000110011011",
    "1110111101101110",
    "1110111001110111",
    "1110111010101111",
    "1110111111011110",
    "1111000110101111",
    "1111001111010010",
    "1111010111111001",
    "1111011111101011",
    "1111100101111110",
    "1111101010011111",
    "1111101101000001",
    "1111101101011101",
    "1111101011100101",
    "1111100111000010",
    "1111011111100011",
    "1111010101000101",
    "1111001000000110",
    "1110111001101101",
    "1110101011100101",
    "1110011111101100",
    "1110011000000100",
    "1110010110011010",
    "1110011011110000",
    "1110101000100101",
    "1110111100011011",
    "1111010101101100",
    "1111110001100101",
    "1111110011011101",
    "1111011101000000",
    "1111001101101110",
    "1111000110110111",
    "1111000111111111",
    "1111001111010100",
    "1111011010010110",
    "1111100110101110",
    "1111110010101111",
    "1111111101100000",
    "1111111001011101",
    "1111110010110000",
    "1111101111000101",
    "1111101111010011",
    "1111110100000011",
    "1111111101011010",
    "1111110101010110",
    "1111100101110111",
    "1111010110000011",
    "1111000111100101",
    "1110111011100101",
    "1110110010010010",
    "1110101011011000",
    "1110100110011011",
    "1110100011001000",
    "1110100001011111",
    "1110100001101001",
    "1110100011110001",
    "1110100111110101",
    "1110101101100000",
    "1110110100001110",
    "1110111011011110",
    "1111000010111011",
    "1111001010110000",
    "1111010011100100",
    "1111011110000000",
    "1111101010100110",
    "1111111001011011",
    "1111110101111110",
    "1111100100100010",
    "1111010011011101",
    "1111000100001000",
    "1110110111110010",
    "1110101111011100",
    "1110101011101000",
    "1110101100011011",
    "1110110001011010",
    "1110111001101111",
    "1111000100010111",
    "1111010000001010",
    "1111011100000100",
    "1111100110111110",
    "1111101111111001",
    "1111110101111000",
    "1111111000001100",
    "1111110110010111",
    "1111110000001111",
    "1111100101111110",
    "1111011000010001",
    "1111001000011101",
    "1110111000011000",
    "1110101010001011",
    "1110011111101011",
    "1110011010001001",
    "1110011001111100",
    "1110011110100011",
    "1110100110111011",
    "1110110001111000",
    "1110111110010100",
    "1111001011010110",
    "1111011000001011",
    "1111100011110110",
    "1111101101010100",
    "1111110011011100",
    "1111110101010001",
    "1111110010011010",
    "1111101011001000",
    "1111100000011100",
    "1111010011111011",
    "1111000111010000",
    "1110111100000001",
    "1110110011010011",
    "1110101101111010",
    "1110101100010001",
    "1110101110101110",
    "1110110101011010",
    "1111000000001101",
    "1111001110101011",
    "1111011111110101",
    "1111110010001111",
    "1111111011110101",
    "1111101100001101",
    "1111100000001111",
    "1111011000100011",
    "1111010101000011",
    "1111010101000110",
    "1111010111110001",
    "1111011100001010",
    "1111100001110000",
    "1111101000000111",
    "1111101111000010",
    "1111110110010000",
    "1111111101010110",
    "1111111100000110",
    "1111110110101000",
    "1111110010011010",
    "1111101111011001",
    "1111101101001101",
    "1111101011010011",
    "1111101001001000",
    "1111100110010101",
    "1111100010110110",
    "1111011110110001",
    "1111011010010011",
    "1111010101101001",
    "1111010000111101",
    "1111001100010100",
    "1111000111111001",
    "1111000011101100",
    "1110111111110011",
    "1110111100010100",
    "1110111001010101",
    "1110110110111100",
    "1110110101011000",
    "1110110100110111",
    "1110110101110001",
    "1110111000010110",
    "1110111101000010",
    "1111000100001010",
    "1111001101111111",
    "1111011010110101",
    "1111101010110010",
    "1111111101011111",
    "1111101110000011",
    "1111011001110101",
    "1111001000010001",
    "1110111011101011",
    "1110110101100111",
    "1110110110010110",
    "1110111100110111",
    "1111000110111111",
    "1111010010011100",
    "1111011101000000",
    "1111100101011101",
    "1111101011000111",
    "1111101101111011",
    "1111101110000010",
    "1111101011101011",
    "1111100111001000",
    "1111100000111000",
    "1111011001101000",
    "1111010010010000",
    "1111001011110011",
    "1111000111000011",
    "1111000100011000",
    "1111000011101001",
    "1111000100010011",
    "1111000101100101",
    "1111000110110100",
    "1111000111011011",
    "1111000111010000",
    "1111000110001110",
    "1111000100100101",
    "1111000010110001",
    "1111000001001111",
    "1111000000100110",
    "1111000001011010",
    "1111000100001011",
    "1111001001001001",
    "1111010000011001",
    "1111011001110000",
    "1111100101000000",
    "1111110001101100",
    "1111111111001111",
    "1111110011001011",
    "1111100110101110",
    "1111011100011011",
    "1111010101000110",
    "1111010001000111",
    "1111010000001010",
    "1111010001010111",
    "1111010011101110",
    "1111010110010011",
    "1111011000110000",
    "1111011011010110",
    "1111011110011110",
    "1111100010100001",
    "1111100111001111",
    "1111101011101100",
    "1111101110011010",
    "1111101101110011",
    "1111101000110111",
    "1111011111101000",
    "1111010011010101",
    "1111000110001101",
    "1110111010101111",
    "1110110011000011",
    "1110110000010101",
    "1110110010110001",
    "1110111001100101",
    "1111000011100010",
    "1111001111011001",
    "1111011100001110",
    "1111101001011111",
    "1111110110111001",
    "1111111011110001",
    "1111101110111101",
    "1111100011010000",
    "1111011001011000",
    "1111010010001010",
    "1111001110001001",
    "1111001101100011",
    "1111010000001111",
    "1111010101110001",
    "1111011101100000",
    "1111100110101111",
    "1111110000101100",
    "1111111010100110",
    "1111111100010010",
    "1111110100110011",
    "1111101111100010",
    "1111101100111001",
    "1111101100111111",
    "1111101111100000",
    "1111110011110011",
    "1111111001000100",
    "1111111110011100",
    "1111111100110011",
    "1111111001001110",
    "1111110111001000",
    "1111110110100110",
    "1111110111100011",
    "1111111001110100",
    "1111111101000110",
    "1111111110111101",
    "1111111010101110",
    "1111110110100000",
    "1111110010100010",
    "1111101110111111",
    "1111101100000010",
    "1111101001111001",
    "1111101000110011",
    "1111101001000111",
    "1111101011000110",
    "1111101110111011",
    "1111110100110001",
    "1111111100100110",
    "1111111001100100",
    "1111101110001001",
    "1111100001110000",
    "1111010101011111",
    "1111001010100110",
    "1111000010011001",
    "1110111101110011",
    "1110111101010010",
    "1111000000111000",
    "1111001000010001",
    "1111010011001101",
    "1111100001001000",
    "1111110000111110",
    "1111111111000011",
    "1111110001010101",
    "1111101000001000",
    "1111100101000110",
    "1111101000101111",
    "1111110010010011",
    "1111111111101110",
    "1111101111001110",
    "1111011101101000",
    "1111001011111010",
    "1110111011000100",
    "1110101100001111",
    "1110100001000101",
    "1110011011010001",
    "1110011100001001",
    "1110100100001011",
    "1110110010100010",
    "1111000101000101",
    "1111011000110111",
    "1111101011000111",
    "1111111001110010",
    "1111111011111010",
    "1111110101110100",
    "1111110010111011",
    "1111110010000100",
    "1111110010010001",
    "1111110011000010",
    "1111110100010100",
    "1111110110010110",
    "1111111001101000",
    "1111111110101001",
    "1111111010000011",
    "1111110000000101",
    "1111100011001101",
    "1111010011101110",
    "1111000010110011",
    "1110110010011001",
    "1110100100100111",
    "1110011011001111",
    "1110010111001000",
    "1110010111110010",
    "1110011011101111",
    "1110100000111001",
    "1110100101100100",
    "1110101000110000",
    "1110101010100101",
    "1110101011110111",
    "1110101101110111",
    "1110110001101011",
    "1110110111110101",
    "1111000000001101",
    "1111001001111101",
    "1111010011110110",
    "1111011100100101",
    "1111100011000000",
    "1111100110010011",
    "1111100101111110",
    "1111100001111110",
    "1111011010110111",
    "1111010001111110",
    "1111001001010011",
    "1111000010111011",
    "1111000000100100",
    "1111000011010101",
    "1111001011010100",
    "1111010111111110",
    "1111101000011000",
    "1111111011100110",
    "1111101111011111",
    "1111011010011110",
    "1111000111010110",
    "1110111000010001",
    "1110101110111111",
    "1110101100010001",
    "1110101111101110",
    "1110110111101111",
    "1111000010000000",
    "1111001100011110",
    "1111010101111110",
    "1111011110100001",
    "1111100111000101",
    "1111110000110111",
    "1111111100101010",
    "1111110101100100",
    "1111100110111001",
    "1111011000110101",
    "1111001101000101",
    "1111000100111011",
    "1111000000111011",
    "1111000001000011",
    "1111000100100010",
    "1111001010010001",
    "1111010000111000",
    "1111010111000011",
    "1111011011100101",
    "1111011101101110",
    "1111011101010010",
    "1111011010100101",
    "1111010110010011",
    "1111010001011100",
    "1111001101000010",
    "1111001010001100",
    "1111001001101111",
    "1111001100010001",
    "1111010010000000",
    "1111011010111000",
    "1111100110100100",
    "1111110100011111",
    "1111111011111011",
    "1111101011011111",
    "1111011011000100",
    "1111001011101000",
    "1110111110010001",
    "1110110011110001",
    "1110101100101010",
    "1110101000111111",
    "1110101000100000",
    "1110101010110010",
    "1110101111100011",
    "1110110110111011",
    "1111000001011001",
    "1111001111010010",
    "1111100000001101",
    "1111110010100100",
    "1111111100000101",
    "1111101110101010",
    "1111100111010111",
    "1111100111001110",
    "1111101101111010",
    "1111111010001111",
    "1111110101000010",
    "1111100000110011",
    "1111001001101101",
    "1110110001000000",
    "1110011000110101",
    "1110000100001101",
    "1101110110000110",
    "1101110000101011",
    "1101110100100101",
    "1110000000111011",
    "1110010011111011",
    "1110101011101111",
    "1111000110101010",
    "1111100011000101",
    "1111111110111110",
    "1111101000010000",
    "1111010101010101",
    "1111001010010011",
    "1111000111110010",
    "1111001100100000",
    "1111010101100101",
    "1111011111100110",
    "1111100111100100",
    "1111101011111110",
    "1111101100110001",
    "1111101011000011",
    "1111101000001100",
    "1111100101000110",
    "1111100001111011",
    "1111011110010110",
    "1111011001110101",
    "1111010100010010",
    "1111001101111010",
    "1111000111010001",
    "1111000001000010",
    "1110111011110000",
    "1110110111111010",
    "1110110101111001",
    "1110110110001001",
    "1110111001001011",
    "1110111111011110",
    "1111001001010101",
    "1111010110101111",
    "1111100111010111",
    "1111111010011101",
    "1111110000101011",
    "1111011010110111",
    "1111000100110001",
    "1110101111000101",
    "1110011010110101",
    "1110001001010000",
    "1101111011100011",
    "1101110010100111",
    "1101101110101000",
    "1101101110111111",
    "1101110010011101",
    "1101110111101101",
    "1101111101101011",
    "1110000100001000",
    "1110001011100011",
    "1110010101001000",
    "1110100010000011",
    "1110110010111001",
    "1111000110111111",
    "1111011100010111",
    "1111110000010001",
    "1111111111101011",
    "1111110111100011",
    "1111110110010111",
    "1111111100000011",
    "1111111001001101",
    "1111101011110011",
    "1111011101111111",
    "1111010001100111",
    "1111001000001011",
    "1111000010101011",
    "1111000001110001",
    "1111000101110100",
    "1111001110011111",
    "1111011010110101",
    "1111101001001001",
    "1111110111010001",
    "1111111100101110",
    "1111110100010010",
    "1111101111110100",
    "1111101110110111",
    "1111110000100100",
    "1111110100000100",
    "1111111001000001",
    "1111111111100100",
    "1111110111101011",
    "1111101100100000",
    "1111011111001111",
    "1111010001001000",
    "1111000100000000",
    "1110111001110100",
    "1110110100010010",
    "1110110100100101",
    "1110111011001110",
    "1111000111111111",
    "1111011010001001",
    "1111110000000110",
    "1111111000011111",
    "1111100010011111",
    "1111010000101011",
    "1111000101001101",
    "1111000001000000",
    "1111000011111000",
    "1111001100100001",
    "1111011001010110",
    "1111101000110010",
    "1111111001110010",
    "1111110100001010",
    "1111100001010100",
    "1111001101111111",
    "1110111011001001",
    "1110101010010001",
    "1110011101000100",
    "1110010100111011",
    "1110010010011010",
    "1110010101001011",
    "1110011100001010",
    "1110100110000100",
    "1110110010000000",
    "1110111111100110",
    "1111001110111111",
    "1111100000001111",
    "1111110010111000",
    "1111111010011001",
    "1111101001110010",
    "1111011101101000",
    "1111010111110010",
    "1111011001000110",
    "1111100001001111",
    "1111101110110110",
    "1111111111111011",
    "1111101101010110",
    "1111011011100101",
    "1111001100110010",
    "1111000010111001",
    "1110111111011010",
    "1111000011000011",
    "1111001101100000",
    "1111011101011100",
    "1111110000110111",
    "1111111010110001",
    "1111101000001111",
    "1111011010000001",
    "1111010010010101",
    "1111010010100111",
    "1111011011010110",
    "1111101011110001",
    "1111111110001100",
    "1111100101101111",
    "1111001110010110",
    "1110111011000111",
    "1110101110000111",
    "1110101000000110",
    "1110101000100010",
    "1110101110001010",
    "1110110111110001",
    "1111000100011010",
    "1111010011101111",
    "1111100101011111",
    "1111111001000111",
    "1111110010010010",
    "1111011110010001",
    "1111001100011011",
    "1110111110001101",
    "1110110100101001",
    "1110110000000101",
    "1110110000010101",
    "1110110100110100",
    "1110111100100101",
    "1111000110101010",
    "1111010001111110",
    "1111011101100000",
    "1111101000010001",
    "1111110001100000",
    "1111111000110000",
    "1111111101111011",
    "1111111110101000",
    "1111111100011111",
    "1111111011000001",
    "1111111001110000",
    "1111111000010001",
    "1111110110010001",
    "1111110011011101",
    "1111101111101101",
    "1111101011000000",
    "1111100101100111",
    "1111100000000111",
    "1111011011010100",
    "1111011000000110",
    "1111010111001001",
    "1111011000111100",
    "1111011101100110",
    "1111100101000101",
    "1111101111001011",
    "1111111011100110",
    "1111110110001000",
    "1111100111000001",
    "1111011000010110",
    "1111001011101011",
    "1111000010001010",
    "1110111100010110",
    "1110111001101101",
    "1110111000111100",
    "1110111000001110",
    "1110110110000011",
    "1110110001011111",
    "1110101010101000",
    "1110100010010100",
    "1110011001110111",
    "1110010010100110",
    "1110001101011001",
    "1110001010101011",
    "1110001010010110",
    "1110001100000101",
    "1110001111101011",
    "1110010101000110",
    "1110011100110111",
    "1110100111100101",
    "1110110101110001",
    "1111000111010011",
    "1111011011001100",
    "1111101111100010",
    "1111111101111110",
    "1111101111100111",
    "1111100110100111",
    "1111100011001000",
    "1111100100010010",
    "1111101000100100",
    "1111101110101000",
    "1111110101100111",
    "1111111101011000",
    "1111111001110011",
    "1111101111110011",
    "1111100100110011",
    "1111011001100000",
    "1111001111000100",
    "1111000110101100",
    "1111000001010100",
    "1110111111010100",
    "1111000000011010",
    "1111000011111100",
    "1111001000111010",
    "1111001110011111",
    "1111010100000000",
    "1111011000111110",
    "1111011101001111",
    "1111100000110101",
    "1111100011101110",
    "1111100110000000",
    "1111100111101010",
    "1111101000101001",
    "1111101000110101",
    "1111101000000111",
    "1111100110011101",
    "1111100011111011",
    "1111100000101100",
    "1111011101000111",
    "1111011001100111",
    "1111010110110010",
    "1111010101010011",
    "1111010101101111",
    "1111011000100011",
    "1111011110000010",
    "1111100110001001",
    "1111110000011001",
    "1111111011101010",
    "1111111001100100",
    "1111110001010101",
    "1111101101100001",
    "1111101111101110",
    "1111111000111000",
    "1111110111001000",
    "1111100001110000",
    "1111001001010011",
    "1110110000110000",
    "1110011011000010",
    "1110001010011101",
    "1110000000010010",
    "1101111100101110",
    "1101111111000111",
    "1110000110001110",
    "1110010000110001",
    "1110011101100001",
    "1110101011010110",
    "1110111001001100",
    "1111000101111110",
    "1111010000101110",
    "1111011000101111",
    "1111011101110010",
    "1111100000001000",
    "1111100000100011",
    "1111100000000111",
    "1111100000000010",
    "1111100001001111",
    "1111100100010000",
    "1111101001000111",
    "1111101111100000",
    "1111110110110010",
    "1111111110001101",
    "1111111011000010",
    "1111110101110101",
    "1111110010101111",
    "1111110010000110",
    "1111110011110111",
    "1111110111101011",
    "1111111100110110",
    "1111111101011001",
    "1111110111111100",
    "1111110011011001",
    "1111110000001000",
    "1111101110010001",
    "1111101101110011",
    "1111101110100111",
    "1111110000101010",
    "1111110011111100",
    "1111111000100000",
    "1111111110010010",
    "1111111010111000",
    "1111110011100110",
    "1111101100100110",
    "1111100110110101",
    "1111100011011010",
    "1111100011010010",
    "1111100110111010",
    "1111101101111001",
    "1111110110111110",
    "1111111111110000",
    "1111111000011001",
    "1111110100101001",
    "1111110101011001",
    "1111111010110001",
    "1111111011011101",
    "1111101101100100",
    "1111011011101101",
    "1111000110101100",
    "1110110000001111",
    "1110011010111111",
    "1110001001111010",
    "1101111111011001",
    "1101111100100011",
    "1110000000101011",
    "1110001001011000",
    "1110010011101001",
    "1110011100110101",
    "1110100100000001",
    "1110101010010100",
    "1110110010010101",
    "1110111110101101",
    "1111010000100011",
    "1111100110101011",
    "1111111101110110",
    "1111101110001011",
    "1111100001001101",
    "1111011101000100",
    "1111100001001000",
    "1111101010110110",
    "1111110111000001",
    "1111111101010001",
    "1111110100000000",
    "1111101110000100",
    "1111101011100001",
    "1111101011111010",
    "1111101110101010",
    "1111110011010110",
    "1111111001100011",
    "1111111111001110",
    "1111110111111010",
    "1111110001011101",
    "1111101100110000",
    "1111101010010111",
    "1111101010011000",
    "1111101100011100",
    "1111110000000001",
    "1111110100011011",
    "1111111000111001",
    "1111111100110000",
    "1111111111011010",
    "1111111111011011",
    "1111111111110000",
    "1111111110110010",
    "1111111100110101",
    "1111111010111110",
    "1111111001100110",
    "1111111000110011",
    "1111111000011101",
    "1111111000010010",
    "1111111000000101",
    "1111110111110010",
    "1111110111100101",
    "1111110111111001",
    "1111111001001111",
    "1111111100001010",
    "1111111110111110",
    "1111110111111011",
    "1111101110010101",
    "1111100001110110",
    "1111010010010101",
    "1111000000001100",
    "1110101100101011",
    "1110011001101010",
    "1110001001100000",
    "1101111110010100",
    "1101111001011110",
    "1101111011011011",
    "1110000011101110",
    "1110010001100010",
    "1110100011111110",
    "1110111010000110",
    "1111010010101100",
    "1111101011110100",
    "1111111101000100",
    "1111101010110011",
    "1111011111011010",
    "1111011011101111",
    "1111011110110011",
    "1111100110010101",
    "1111101111011110",
    "1111110111101100",
    "1111111101100011",
    "1111111111010000",
    "1111111110010010",
    "1111111110101001",
    "1111111111100100",
    "1111111111011011",
    "1111111110101111",
    "1111111110101001",
    "1111111111011101",
    "1111111110100010",
    "1111111011001111",
    "1111110110111001",
    "1111110010000011",
    "1111101101011101",
    "1111101001110000",
    "1111100111001101",
    "1111100101101100",
    "1111100100110011",
    "1111100011111100",
    "1111100010100110",
    "1111100000010010",
    "1111011100110000",
    "1111010111110100",
    "1111010001010000",
    "1111001000111111",
    "1110111110111111",
    "1110110011100010",
    "1110100111010110",
    "1110011011101000",
    "1110010001100110",
    "1110001010011011",
    "1110000110101010",
    "1110000110010000",
    "1110001000100111",
    "1110001100111000",
    "1110010010010000",
    "1110011000010101",
    "1110011111000111",
    "1110100111101010",
    "1110110011101010",
    "1111000100110111",
    "1111011011101111",
    "1111110110110111",
    "1111101101000111",
    "1111010100110110",
    "1111000100100010",
    "1110111110111010",
    "1111000100000110",
    "1111010001111101",
    "1111100101011000",
    "1111111011011010",
    "1111101110000100",
    "1111011000101100",
    "1111000101101110",
    "1110110110100101",
    "1110101100110010",
    "1110101001011110",
    "1110101101000010",
    "1110110110101100",
    "1111000100101100",
    "1111010100111001",
    "1111100101011000",
    "1111110100111110",
    "1111111100111001",
    "1111110000101011",
    "1111100110111101",
    "1111100000110000",
    "1111011111000000",
    "1111100010010000",
    "1111101001111101",
    "1111110100101010",
    "1111111111100111",
    "1111110101000100",
    "1111101101001010",
    "1111101000110001",
    "1111101000010000",
    "1111101011110110",
    "1111110011111010",
    "1111111111011001",
    "1111101110100101",
    "1111011010111111",
    "1111000110101101",
    "1110110100010101",
    "1110100110000100",
    "1110011101011100",
    "1110011010101111",
    "1110011101001111",
    "1110100011101110",
    "1110101100111100",
    "1110110111111111",
    "1111000100010111",
    "1111010001100010",
    "1111011110111010",
    "1111101011101000",
    "1111110110110011",
    "1111111111100111",
    "1111111010010001",
    "1111110111000011",
    "1111110110011110",
    "1111111000011100",
    "1111111101001011",
    "1111111010111000",
    "1111101111100011",
    "1111100001000111",
    "1111010000100111",
    "1110111111111000",
    "1110110000110110",
    "1110100101001110",
    "1110011110000010",
    "1110011011011011",
    "1110011100110010",
    "1110100001001111",
    "1110101000000011",
    "1110110001000111",
    "1110111100110111",
    "1111001011101101",
    "1111011101100001",
    "1111110001000010",
    "1111111100000000",
    "1111101100101111",
    "1111100011111011",
    "1111100011010101",
    "1111101011000010",
    "1111111001100010",
    "1111110011101111",
    "1111100000001000",
    "1111001110110011",
    "1111000010010101",
    "1110111100011011",
    "1110111101100110",
    "1111000101011101",
    "1111010010111001",
    "1111100100010111",
    "1111110111111101",
    "1111110100001101",
    "1111100010001000",
    "1111010011010101",
    "1111001000111110",
    "1111000011100001",
    "1111000010101110",
    "1111000101101100",
    "1111001011001111",
    "1111010010000101",
    "1111011001010001",
    "1111100000010001",
    "1111100111000101",
    "1111101110000010",
    "1111110101101110",
    "1111111110101010",
    "1111110110110010",
    "1111101010111000",
    "1111011110010010",
    "1111010010010010",
    "1111001000011011",
    "1111000010010101",
    "1111000001001000",
    "1111000101010010",
    "1111001110011001",
    "1111011011010001",
    "1111101010011010",
    "1111111010011011",
    "1111110101100111",
    "1111100110011010",
    "1111011000011101",
    "1111001100011011",
    "1111000011000011",
    "1110111101000100",
    "1110111010110100",
    "1110111100000001",
    "1110111111111101",
    "1111000101100101",
    "1111001011111101",
    "1111010010101011",
    "1111011001110100",
    "1111100001111011",
    "1111101011100000",
    "1111110110100101",
    "1111111101100110",
    "1111110010101011",
    "1111101010110010",
    "1111100111111100",
    "1111101011011110",
    "1111110101011010",
    "1111111011101000",
    "1111101010011100",
    "1111011010001111",
    "1111001110001010",
    "1111001000011000",
    "1111001001110101",
    "1111010010000010",
    "1111011111100011",
    "1111110000011011",
    "1111111101010101",
    "1111101011101111",
    "1111011100100000",
    "1111010001001101",
    "1111001011001010",
    "1111001011001110",
    "1111010001100110",
    "1111011101100011",
    "1111101101010111",
    "1111111110100110",
    "1111110001011000",
    "1111100100110011",
    "1111011100110010",
    "1111011001011000",
    "1111011001100101",
    "1111011011111100",
    "1111011111010010",
    "1111100011010010",
    "1111101000101001",
    "1111110000111000",
    "1111111101011100",
    "1111110001000000",
    "1111011011011000",
    "1111000011111001",
    "1110101101110111",
    "1110011100101101",
    "1110010011000001",
    "1110010001111101",
    "1110011000111010",
    "1110100110000100",
    "1110110110111110",
    "1111001001000100",
    "1111011010010001",
    "1111101001001000",
    "1111110100110011",
    "1111111100111110",
    "1111111110010000",
    "1111111100101110",
    "1111111110000011",
    "1111111110001101",
    "1111111000100101",
    "1111110001011011",
    "1111101001000110",
    "1111011111111011",
    "1111010110010010",
    "1111001100101011",
    "1111000011101100",
    "1110111011111010",
    "1110110101101100",
    "1110110001010000",
    "1110101110101000",
    "1110101101101101",
    "1110101110101001",
    "1110110001110011",
    "1110110111111110",
    "1111000010000010",
    "1111010000100100",
    "1111100011001101",
    "1111111000001110",
    "1111110011010110",
    "1111100011000110",
    "1111011010000010",
    "1111011001110010",
    "1111100010000010",
    "1111110000110111",
    "1111111100100100",
    "1111101001011000",
    "1111011000001000",
    "1111001010110101",
    "1111000011001010",
    "1111000010001000",
    "1111001000001100",
    "1111010100111011",
    "1111100110101110",
    "1111111011000111",
    "1111110000111000",
    "1111100000001010",
    "1111010100100010",
    "1111001110100001",
    "1111001101011110",
    "1111010000000010",
    "1111010100110110",
    "1111011011000010",
    "1111100010011111",
    "1111101011011111",
    "1111110110011110",
    "1111111100010110",
    "1111101101010001",
    "1111011100111100",
    "1111001100011011",
    "1110111100110111",
    "1110101111001111",
    "1110100100010111",
    "1110011100101010",
    "1110011000001110",
    "1110010110110111",
    "1110011000001011",
    "1110011011101011",
    "1110100000111000",
    "1110100111010000",
    "1110101110011011",
    "1110110110001001",
    "1110111110011110",
    "1111000111100010",
    "1111010001100100",
    "1111011100101101",
    "1111101001000000",
    "1111110110010110",
    "1111111011100000",
    "1111101101010000",
    "1111011111110001",
    "1111010100001011",
    "1111001011011000",
    "1111000110000011",
    "1111000100001110",
    "1111000101011111",
    "1111001000111010",
    "1111001101011100",
    "1111010010000110",
    "1111010110001000",
    "1111011000110111",
    "1111011001101011",
    "1111011000000100",
    "1111010011101001",
    "1111001100100000",
    "1111000011011000",
    "1110111001101101",
    "1110110001010010",
    "1110101011111010",
    "1110101010110111",
    "1110101110101101",
    "1110110111001001",
    "1111000011100010",
    "1111010011000000",
    "1111100100110001",
    "1111110111110101",
    "1111110101001010",
    "1111100100000001",
    "1111010110100101",
    "1111001110001010",
    "1111001011001110",
    "1111001101001010",
    "1111010010011100",
    "1111011001010001",
    "1111100000001000",
    "1111100110010000",
    "1111101011100010",
    "1111110000001010",
    "1111110100001101",
    "1111110111010000",
    "1111111000100101",
    "1111110111010001",
    "1111110010110101",
    "1111101011010101",
    "1111100001101001",
    "1111010111000011",
    "1111001100111010",
    "1111000100010101",
    "1110111101110101",
    "1110111001100101",
    "1110110111011111",
    "1110110111010101",
    "1110111000111100",
    "1110111100001100",
    "1111000000111000",
    "1111000110101100",
    "1111001101001010",
    "1111010011111000",
    "1111011010011000",
    "1111100000100100",
    "1111100110011100",
    "1111101100010011",
    "1111110010100000",
    "1111111001010111",
    "1111111110111001",
    "1111110110010100",
    "1111101101000001",
    "1111100011010111",
    "1111011001111001",
    "1111010001011010",
    "1111001010110111",
    "1111000110110111",
    "1111000101101100",
    "1111000110110111",
    "1111001001010011",
    "1111001011010011",
    "1111001011000110",
    "1111000111001101",
    "1110111110110101",
    "1110110010001000",
    "1110100010011100",
    "1110010001110100",
    "1110000010110100",
    "1101110111110010",
    "1101110010011001",
    "1101110011011101",
    "1101111011000100",
    "1110001000101100",
    "1110011011011101",
    "1110110010000101",
    "1111001010111010",
    "1111100011101001",
    "1111111001100010",
    "1111110101111011",
    "1111101100101011",
    "1111101011001010",
    "1111110000010111",
    "1111111010000010",
    "1111111010100011",
    "1111110000000110",
    "1111101000010011",
    "1111100011111100",
    "1111100010111000",
    "1111100100010011",
    "1111100111010111",
    "1111101011001010",
    "1111101111000101",
    "1111110010101110",
    "1111110101110100",
    "1111111000001010",
    "1111111001101101",
    "1111111010011101",
    "1111111010100001",
    "1111111001111001",
    "1111111000100011",
    "1111110110010000",
    "1111110010101010",
    "1111101101011010",
    "1111100110011000",
    "1111011101110010",
    "1111010100001011",
    "1111001010010110",
    "1111000001001010",
    "1110111001010000",
    "1110110010110110",
    "1110101101111011",
    "1110101010001100",
    "1110100111010110",
    "1110100101001001",
    "1110100011100100",
    "1110100010100001",
    "1110100010000011",
    "1110100010000000",
    "1110100010010010",
    "1110100010111001",
    "1110100100000110",
    "1110100110100100",
    "1110101011001001",
    "1110110010110011",
    "1110111101111111",
    "1111001100010100",
    "1111011100010100",
    "1111101011100110",
    "1111110111101011",
    "1111111110100110",
    "1111111111101110",
    "1111111011110001",
    "1111110100011011",
    "1111101011101100",
    "1111100011000101",
    "1111011011001100",
    "1111010100000000",
    "1111001101010010",
    "1111000111011000",
    "1111000011001111",
    "1111000010001000",
    "1111000101001110",
    "1111001100111100",
    "1111011000110100",
    "1111100111101001",
    "1111111000000000",
    "1111110111100010",
    "1111101000001011",
    "1111011010110000",
    "1111001111111111",
    "1111001000011101",
    "1111000100101100",
    "1111000101000001",
    "1111001001100111",
    "1111010010010000",
    "1111011110110000",
    "1111101110011101",
    "1111111111100110",
    "1111101100111100",
    "1111011011010011",
    "1111001100010100",
    "1111000001010100",
    "1110111010110100",
    "1110111000100101",
    "1110111001100111",
    "1110111100100011",
    "1111000000001000",
    "1111000011100010",
    "1111000110011010",
    "1111001000111001",
    "1111001011010011",
    "1111001101111111",
    "1111010001010100",
    "1111010101011101",
    "1111011010100101",
    "1111100000100110",
    "1111100111010101",
    "1111101110001110",
    "1111110100100011",
    "1111111001100000",
    "1111111100011111",
    "1111111101010100",
    "1111111100011100",
    "1111111010101111",
    "1111111001010110",
    "1111111001011000",
    "1111111011101110",
    "1111111111001001",
    "1111110111001111",
    "1111101100110001",
    "1111100000001100",
    "1111010010001101",
    "1111000011111110",
    "1110110111001000",
    "1110101101101011",
    "1110101001110100",
    "1110101101010010",
    "1110111001000110",
    "1111001100100001",
    "1111100101001011",
    "1111111111010010",
    "1111101001001001",
    "1111010111100010",
    "1111001101101000",
    "1111001011010110",
    "1111001110111011",
    "1111010101110110",
    "1111011101101101",
    "1111100101010101",
    "1111101100111101",
    "1111110101101010",
    "1111111111010111",
    "1111110001101110",
    "1111100010000000",
    "1111010001110000",
    "1111000010111001",
    "1110110110111111",
    "1110101110101101",
    "1110101001101000",
    "1110100110100100",
    "1110100100000110",
    "1110100001001100",
    "1110011101010010",
    "1110011000011101",
    "1110010011000000",
    "1110001101101000",
    "1110001000110101",
    "1110000101000101",
    "1110000010011101",
    "1110000001000010",
    "1110000000101100",
    "1110000001010010",
    "1110000010100100",
    "1110000100001011",
    "1110000101110110",
    "1110000111100000",
    "1110001001001001",
    "1110001011000010",
    "1110001101010111",
    "1110010000011110",
    "1110010100100000",
    "1110011001101010",
    "1110100000001010",
    "1110101000010110",
    "1110110010101100",
    "1110111111101001",
    "1111001111010010",
    "1111100000111011",
    "1111110011000010",
    "1111111100011111",
    "1111101111110111",
    "1111101000100101",
    "1111100111000101",
    "1111101010101001",
    "1111110001110010",
    "1111111011000001",
    "1111111010011110",
    "1111101110101000",
    "1111100000100110",
    "1111001111110110",
    "1110111101000101",
    "1110101010100011",
    "1110011011011001",
    "1110010010101011",
    "1110010010001000",
    "1110011001101011",
    "1110100111110001",
    "1110111010000100",
    "1111001110110000",
    "1111100100110110",
    "1111111011101011",
    "1111101101101100",
    "1111011001000111",
    "1111001000111001",
    "1110111111000100",
    "1110111100100110",
    "1111000001000010",
    "1111001010011000",
    "1111010110000100",
    "1111100001111110",
    "1111101100111001",
    "1111110110111010",
    "1111111111010001",
    "1111110101001101",
    "1111101011000111",
    "1111100010001010",
    "1111011011110111",
    "1111011001100000",
    "1111011011010100",
    "1111100000011001",
    "1111100110111000",
    "1111101100100110",
    "1111101111100111",
    "1111101110101101",
    "1111101001100011",
    "1111100000100100",
    "1111010100101111",
    "1111000111010110",
    "1110111001101011",
    "1110101100110111",
    "1110100001110011",
    "1110011001000110",
    "1110010011001111",
    "1110010000011110",
    "1110010000111101",
    "1110010100101010",
    "1110011011011110",
    "1110100101001101",
    "1110110001101100",
    "1111000000101011",
    "1111010001101100",
    "1111100100001010",
    "1111110111010001",
    "1111110101100111",
    "1111100011010000",
    "1111010010001010",
    "1111000011000000",
    "1110110110100000",
    "1110101101100110",
    "1110101001000010",
    "1110101001010011",
    "1110101110011100",
    "1110111000001011",
    "1111000101110100",
    "1111010110010011",
    "1111101000001010",
    "1111111001011101",
    "1111111000000110",
    "1111101110111011",
    "1111101101000111",
    "1111110011111100",
    "1111111100101110",
    "1111100110111010",
    "1111001101111111",
    "1110110110000001",
    "1110100010101001",
    "1110010110010000",
    "1110010001100010",
    "1110010011100100",
    "1110011010101010",
    "1110100101011111",
    "1110110011110110",
    "1111000110000001",
    "1111011011110111",
    "1111110011111110",
    "1111110100100000",
    "1111100001010111",
    "1111010110000110",
    "1111010100110100",
    "1111011101011100",
    "1111101101110111",
    "1111111101001100",
    "1111100111010001",
    "1111010011010000",
    "1111000011000101",
    "1110110111110101",
    "1110110001111011",
    "1110110001100001",
    "1110110110011010",
    "1111000000001100",
    "1111001110000000",
    "1111011110110000",
    "1111110001000001",
    "1111111100100111",
    "1111101011011100",
    "1111011100010011",
    "1111001111110011",
    "1111000110011010",
    "1111000000011001",
    "1110111101111000",
    "1110111110100110",
    "1111000010000011",
    "1111000111100000",
    "1111001110001111",
    "1111010101101100",
    "1111011101100011",
    "1111100101101100",
    "1111101110010100",
    "1111110111101101",
    "1111111101110010",
    "1111110001111110",
    "1111100100101001",
    "1111010101101110",
    "1111000101100100",
    "1110110100111110",
    "1110100101011000",
    "1110011000011011",
    "1110001111100001",
    "1110001011011011",
    "1110001100001001",
    "1110010001000010",
    "1110011001000110",
    "1110100011101010",
    "1110110000100011",
    "1110111111110110",
    "1111010001010111",
    "1111100100001000",
    "1111110110001001",
    "1111111010111010",
    "1111110001001101",
    "1111101101110111",
    "1111110000100101",
    "1111110111110100",
    "1111111110101010",
    "1111110101010000",
    "1111101101110000",
    "1111101001010101",
    "1111101000011111",
    "1111101011001111",
    "1111110001001101",
    "1111111001101011",
    "1111111100011001",
    "1111110010011100",
    "1111101001110000",
    "1111100011010101",
    "1111011111101000",
    "1111011110100011",
    "1111011111100110",
    "1111100010010000",
    "1111100110001110",
    "1111101011101011",
    "1111110010111000",
    "1111111100000101",
    "1111111000111001",
    "1111101100111110",
    "1111100001011110",
    "1111011000000001",
    "1111010010001101",
    "1111010001001000",
    "1111010101010000",
    "1111011110000111",
    "1111101010100011",
    "1111111000111110",
    "1111111000011000",
    "1111101011001010",
    "1111100000100100",
    "1111011001011000",
    "1111010101110100",
    "1111010101110010",
    "1111011000111100",
    "1111011110110001",
    "1111100110110010",
    "1111110000011110",
    "1111111011011101",
    "1111111000100010",
    "1111101011110011",
    "1111011110100100",
    "1111010001001100",
    "1111000100001011",
    "1110111000001100",
    "1110101101111011",
    "1110100110000000",
    "1110100000110101",
    "1110011110101000",
    "1110011111010111",
    "1110100010111001",
    "1110101000111001",
    "1110110001000011",
    "1110111010110111",
    "1111000101100101",
    "1111010000000010",
    "1111011000101111",
    "1111011110000101",
    "1111011110101011",
    "1111011001110000",
    "1111001111101001",
    "1111000001111101",
    "1110110011010011",
    "1110100110110110",
    "1110011111010100",
    "1110011110101001",
    "1110100101101010",
    "1110110100010011",
    "1111001001111001",
    "1111100101010101",
    "1111111011001111",
    "1111011010101111",
    "1110111100110010",
    "1110100101000101",
    "1110010110100100",
    "1110010010011001",
    "1110010111101101",
    "1110100011111001",
    "1110110011101100",
    "1111000100000101",
    "1111010011001000",
    "1111100000000101",
    "1111101010111110",
    "1111110100000110",
    "1111111011101100",
    "1111111110010101",
    "1111111010010100",
    "1111111000001111",
    "1111110111101010",
    "1111110111101011",
    "1111110111001000",
    "1111110101000100",
    "1111110001001100",
    "1111101011111001",
    "1111100110001011",
    "1111100001000101",
    "1111011101011001",
    "1111011011011011",
    "1111011011000001",
    "1111011011101011",
    "1111011101000111",
    "1111011111001101",
    "1111100010011100",
    "1111100111011011",
    "1111101110110100",
    "1111111000101001",
    "1111111011110001",
    "1111101111111110",
    "1111100101101100",
    "1111011110011111",
    "1111011011010100",
    "1111011100010100",
    "1111100000111001",
    "1111100111111110",
    "1111110000010001",
    "1111111000011101",
    "1111111111010010",
    "1111111100010011",
    "1111111011001010",
    "1111111101101000",
    "1111111100011110",
    "1111110100000011",
    "1111101010011011",
    "1111100001001000",
    "1111011001100101",
    "1111010100101111",
    "1111010011000101",
    "1111010100011010",
    "1111011000010101",
    "1111011110001101",
    "1111100101011010",
    "1111101101010010",
    "1111110101000001",
    "1111111011101110",
    "1111111111101000",
    "1111111110000101",
    "1111111111101101",
    "1111111001101100",
    "1111110000011001",
    "1111100100111100",
    "1111011000110010",
    "1111001101010110",
    "1111000011101001",
    "1110111100001111",
    "1110110111010011",
    "1110110100110100",
    "1110110100101111",
    "1110110111010001",
    "1110111100111010",
    "1111000110000100",
    "1111010010111110",
    "1111100011001111",
    "1111110101101010",
    "1111110111100010",
    "1111100110011011",
    "1111011000110010",
    "1111001111101110",
    "1111001011011101",
    "1111001011011011",
    "1111001110100011",
    "1111010011100010",
    "1111011001010001",
    "1111011110101101",
    "1111100011000011",
    "1111100101101111",
    "1111100110011101",
    "1111100101001001",
    "1111100010001101",
    "1111011110001010",
    "1111011001110101",
    "1111010101111001",
    "1111010011000011",
    "1111010001101001",
    "1111010001111001",
    "1111010011110001",
    "1111010111000011",
    "1111011011011110",
    "1111100000101100",
    "1111100110010101",
    "1111101011111110",
    "1111110001010111",
    "1111110110011101",
    "1111111011100000",
    "1111111111000001",
    "1111111000110010",
    "1111110001100110",
    "1111101001101111",
    "1111100010000010",
    "1111011011101000",
    "1111010111110001",
    "1111010111011101",
    "1111011011001010",
    "1111100010111001",
    "1111101110010100",
    "1111111100111010",
    "1111110010000001",
    "1111011111100110",
    "1111001101011110",
    "1110111101110000",
    "1110110010100110",
    "1110101101100100",
    "1110101111000111",
    "1110110110010011",
    "1111000001001100",
    "1111001101001110",
    "1111011000010000",
    "1111100000110001",
    "1111100110001101",
    "1111101000101101",
    "1111101000101110",
    "1111100110111011",
    "1111100011111011",
    "1111100000010010",
    "1111011100101101",
    "1111011001111010",
    "1111011000110100",
    "1111011010011000",
    "1111011111011001",
    "1111101000010110",
    "1111110101001011",
    "1111111010101101",
    "1111101000101110",
    "1111010110101101",
    "1111000111000011",
    "1110111011110111",
    "1110110110101111",
    "1110111000000100",
    "1110111111001010",
    "1111001010001011",
    "1111010110110010",
    "1111100010100111",
    "1111101011110010",
    "1111110001010010",
    "1111110010111000",
    "1111110001000000",
    "1111101100011000",
    "1111100101111100",
    "1111011110100100",
    "1111010111001110",
    "1111010000111101",
    "1111001100111101",
    "1111001100010011",
    "1111001111100011",
    "1111010110101100",
    "1111100000110001",
    "1111101100010001",
    "1111110111100010",
    "1111111110110101",
    "1111110111101011",
    "1111110011000011",
    "1111110000100100",
    "1111101111100110",
    "1111101111110001",
    "1111110001010000",
    "1111110100111011",
    "1111111100000011",
    "1111111000010011",
    "1111101000000010",
    "1111010100011101",
    "1111000000010101",
    "1110101111001100",
    "1110100100010101",
    "1110100001101100",
    "1110100111011111",
    "1110110100001110",
    "1111000101010111",
    "1111011000000100",
    "1111101001110110",
    "1111111000111011",
    "1111111011111011",
    "1111110101100100",
    "1111110100010111",
    "1111111000011111",
    "1111111110010001",
    "1111110000101111",
    "1111100000000011",
    "1111001101111000",
    "1110111011110111",
    "1110101011100001",
    "1110011110000000",
    "1110010011111001",
    "1110001101010110",
    "1110001010001011",
    "1110001001111100",
    "1110001100001100",
    "1110010000010111",
    "1110010101110110",
    "1110011100001001",
    "1110100010110110",
    "1110101001100111",
    "1110110000001100",
    "1110110110010101",
    "1110111011101111",
    "1111000000000101",
    "1111000011001111",
    "1111000101000101",
    "1111000101110110",
    "1111000101111100",
    "1111000110000011",
    "1111000110110001",
    "1111001000101000",
    "1111001011111000",
    "1111010000011001",
    "1111010101111001",
    "1111011011111101",
    "1111100010010111",
    "1111101000111010",
    "1111101111100000",
    "1111110101111011",
    "1111111011111001",
    "1111111111000001",
    "1111111011010010",
    "1111111001000100",
    "1111111000010010",
    "1111111000101101",
    "1111111010000010",
    "1111111100001011",
    "1111111111010101",
    "1111111100000011",
    "1111110101101011",
    "1111101101011100",
    "1111100011111001",
    "1111011010001001",
    "1111010001101011",
    "1111001011110111",
    "1111001001111001",
    "1111001100010011",
    "1111010011010010",
    "1111011110110000",
    "1111101110011110",
    "1111111110001101",
    "1111101000110011",
    "1111010011011100",
    "1111000000101110",
    "1110110011000110",
    "1110101100001110",
    "1110101100011011",
    "1110110010110100",
    "1110111101011011",
    "1111001010000010",
    "1111010110101000",
    "1111100001100010",
    "1111101001101000",
    "1111101110000011",
    "1111101110011100",
    "1111101010110110",
    "1111100011111110",
    "1111011011001110",
    "1111010010100110",
    "1111001100001111",
    "1111001001111101",
    "1111001100101011",
    "1111010100001010",
    "1111011111000111",
    "1111101011101010",
    "1111110111110110",
    "1111111101110011",
    "1111110110001101",
    "1111110001011010",
    "1111101110110111",
    "1111101101101110",
    "1111101101000001",
    "1111101011111111",
    "1111101010000101",
    "1111100111000101",
    "1111100011000101",
    "1111011110011100",
    "1111011001110111",
    "1111010110000001",
    "1111010011100111",
    "1111010011001101",
    "1111010101000101",
    "1111011001001100",
    "1111011111011110",
    "1111100111101111",
    "1111110010000101",
    "1111111110101011",
    "1111110010001100",
    "1111100000101011",
    "1111001101011100",
    "1110111010000100",
    "1110101000101000",
    "1110011011011001",
    "1110010011111011",
    "1110010010111011",
    "1110011000010110",
    "1110100011101010",
    "1110110100001011",
    "1111001001001110",
    "1111100001011010",
    "1111111010100000",
    "1111101110100110",
    "1111011101000111",
    "1111010011011000",
    "1111010010000101",
    "1111011000000100",
    "1111100010110100",
    "1111101111011000",
    "1111111011011110",
    "1111111001111110",
    "1111110001001101",
    "1111101001110111",
    "1111100011110001",
    "1111011111010001",
    "1111011101000111",
    "1111011110001101",
    "1111100010110011",
    "1111101010001111",
    "1111110011000110",
    "1111111011100011",
    "1111111101110101",
    "1111111001111011",
    "1111111000100111",
    "1111111001011010",
    "1111111011101110",
    "1111111111001101",
    "1111111100001001",
    "1111110110001111",
    "1111101110110010",
    "1111100101101110",
    "1111011011001100",
    "1111001111111011",
    "1111000100111110",
    "1110111011101000",
    "1110110101001110",
    "1110110010110011",
    "1110110100110110",
    "1110111011000010",
    "1111000100011100",
    "1111001111011010",
    "1111011010000111",
    "1111100010110110",
    "1111101000011000",
    "1111101010010000",
    "1111101000101110",
    "1111100100100100",
    "1111011110101101",
    "1111011000000001",
    "1111010001000101",
    "1111001010001100",
    "1111000011011010",
    "1110111100100110",
    "1110110101100101",
    "1110101110010001",
    "1110100110101010",
    "1110011111000000",
    "1110010111110001",
    "1110010001100110",
    "1110001101001100",
    "1110001011001110",
    "1110001100001100",
    "1110010000011100",
    "1110011000000001",
    "1110100010110001",
    "1110110000001111",
    "1110111111100100",
    "1111001111100011",
    "1111011110011110",
    "1111101010100000",
    "1111110010000000",
    "1111110011110011",
    "1111101111100000",
    "1111100101101111",
    "1111011000001011",
    "1111001001000111",
    "1110111011001110",
    "1110110000110000",
    "1110101011010001",
    "1110101011011001",
    "1110110000111011",
    "1110111011000110",
    "1111001000111001",
    "1111011001001011",
    "1111101010100011",
    "1111111011010101",
    "1111110110010010",
    "1111101100001100",
    "1111100111100000",
    "1111101000100010",
    "1111101110101000",
    "1111111000011000",
    "1111111011110101",
    "1111101111110010",
    "1111100100101111",
    "1111011011110010",
    "1111010101011101",
    "1111010010001010",
    "1111010010000011",
    "1111010101000001",
    "1111011010100110",
    "1111100010001011",
    "1111101010110111",
    "1111110011110110",
    "1111111100100100",
    "1111111011001001",
    "1111110011001000",
    "1111101010111110",
    "1111100010010111",
    "1111011001010101",
    "1111010000001101",
    "1111000111110001",
    "1111000000110000",
    "1110111011110111",
    "1110111001101010",
    "1110111010010001",
    "1110111101101101",
    "1111000011110100",
    "1111001100100001",
    "1111010111111010",
    "1111100110000100",
    "1111110110111010",
    "1111110110010010",
    "1111100011000110",
    "1111010001100110",
    "1111000011101100",
    "1110111010110100",
    "1110110111010011",
    "1110111000100000",
    "1110111101001010",
    "1111000011111110",
    "1111001100001001",
    "1111010101101001",
    "1111100000111110",
    "1111101110110000",
    "1111111110111010",
    "1111101111011101",
    "1111011110011001",
    "1111010000011100",
    "1111000111111110",
    "1111000110011010",
    "1111001011111100",
    "1111010111001110",
    "1111100101111011",
    "1111110101000111",
    "1111111101111000",
    "1111110101010001",
    "1111110010000110",
    "1111110100011001",
    "1111111011001100",
    "1111111011001010",
    "1111110000110000",
    "1111100111011100",
    "1111100000110000",
    "1111011101100011",
    "1111011110001001",
    "1111100010010100",
    "1111101001010111",
    "1111110010011111",
    "1111111100101110",
    "1111111000101101",
    "1111101110100111",
    "1111100101100101",
    "1111011110000010",
    "1111011000001100",
    "1111010100000110",
    "1111010001011111",
    "1111010000000111",
    "1111001111111111",
    "1111010001101011",
    "1111010110001011",
    "1111011110110011",
    "1111101100010111",
    "1111111110111101",
    "1111101010011001",
    "1111010001101110",
    "1110111001101010",
    "1110100100101100",
    "1110010100101010",
    "1110001010011000",
    "1110000101011111",
    "1110000100111001",
    "1110000111001001",
    "1110001010111100",
    "1110001111010110",
    "1110010011110100",
    "1110011000010001",
    "1110011100101110",
    "1110100001001111",
    "1110100101110110",
    "1110101010011110",
    "1110101111001010",
    "1110110011110011",
    "1110111000010000",
    "1110111100010110",
    "1110111111110101",
    "1111000010010100",
    "1111000011011100",
    "1111000011000101",
    "1111000001010101",
    "1110111110110101",
    "1110111100100011",
    "1110111011110011",
    "1110111110000111",
    "1111000100111001",
    "1111010001001100",
    "1111100010111001",
    "1111111000010110",
    "1111110001011111",
    "1111011110011011",
    "1111010001101100",
    "1111001101001100",
    "1111010000110001",
    "1111011010100000",
    "1111100111011001",
    "1111110100101010",
    "1111111111001101",
    "1111110100011111",
    "1111101010011001",
    "1111100000001111",
    "1111010110001000",
    "1111001101001110",
    "1111000111010101",
    "1111000110010000",
    "1111001010110100",
    "1111010100010010",
    "1111100000101001",
    "1111101101010010",
    "1111110111110101",
    "1111111110111101",
    "1111111101101000",
    "1111111101011111",
    "1111111111111001",
    "1111111011110001",
    "1111110101111111",
    "1111101111000001",
    "1111100111001011",
    "1111011111000000",
    "1111010111010011",
    "1111010000101100",
    "1111001011101101",
    "1111001000010000",
    "1111000101111100",
    "1111000100001110",
    "1111000010101001",
    "1111000000111001",
    "1110111110110110",
    "1110111100011110",
    "1110111001110100",
    "1110110110110111",
    "1110110011101110",
    "1110110000101100",
    "1110101110001101",
    "1110101100110010",
    "1110101100110010",
    "1110101110010001",
    "1110110001001000",
    "1110110101001000",
    "1110111010001001",
    "1111000000001010",
    "1111000111010001",
    "1111001111100100",
    "1111011000110100",
    "1111100010011111",
    "1111101011110110",
    "1111110100000101",
    "1111111010101100",
    "1111111111100010",
    "1111111100111101",
    "1111111010001001",
    "1111110111001100",
    "1111110011010010",
    "1111101101110001",
    "1111100110010010",
    "1111011100101110",
    "1111010001100010",
    "1111000101100111",
    "1110111010000111",
    "1110110000011010",
    "1110101001101011",
    "1110100110100100",
    "1110100111000001",
    "1110101010100010",
    "1110110000001010",
    "1110110110111110",
    "1110111110001111",
    "1111000101100000",
    "1111001100101010",
    "1111010011101110",
    "1111011010110111",
    "1111100010000110",
    "1111101001011111",
    "1111110000111001",
    "1111111000001010",
    "1111111111000111",
    "1111111010011010",
    "1111110100110000",
    "1111110000000110",
    "1111101100100110",
    "1111101010011011",
    "1111101001101010",
    "1111101010010110",
    "1111101100011100",
    "1111101111110111",
    "1111110100011100",
    "1111111001111001",
    "1111111111111101",
    "1111111001101001",
    "1111110011010001",
    "1111101101001010",
    "1111100111100100",
    "1111100010101110",
    "1111011110111000",
    "1111011100001110",
    "1111011010111100",
    "1111011011010011",
    "1111011101010110",
    "1111100001001101",
    "1111100110101011",
    "1111101101011001",
    "1111110100101001",
    "1111111011100000",
    "1111111110111011",
    "1111111011100001",
    "1111111010101010",
    "1111111100001110",
    "1111111111100101",
    "1111111100001111",
    "1111111000100011",
    "1111110110011000",
    "1111110110100000",
    "1111111001000110",
    "1111111101110011",
    "1111111100001011",
    "1111110110000011",
    "1111110000111001",
    "1111101101101000",
    "1111101100111001",
    "1111101110111110",
    "1111110011111101",
    "1111111011110010",
    "1111111001100011",
    "1111101100010110",
    "1111011101001010",
    "1111001101010001",
    "1110111110101110",
    "1110110011110100",
    "1110101110101000",
    "1110110000011111",
    "1110111001101000",
    "1111001001000001",
    "1111011100101010",
    "1111110001110111",
    "1111111010000000",
    "1111101001010001",
    "1111011101001111",
    "1111010110010011",
    "1111010011110110",
    "1111010100100000",
    "1111010110100101",
    "1111011000011010",
    "1111011000101111",
    "1111010110111111",
    "1111010011010011",
    "1111001110010001",
    "1111001000111001",
    "1111000100001000",
    "1111000000110001",
    "1110111111001000",
    "1110111111001111",
    "1111000000110001",
    "1111000011010111",
    "1111000110101101",
    "1111001010100110",
    "1111001110111010",
    "1111010011100110",
    "1111011000101010",
    "1111011110000111",
    "1111100011111011",
    "1111101001111000",
    "1111101111110101",
    "1111110101101000",
    "1111111011001101",
    "1111111111010011",
    "1111111001111010",
    "1111110100011000",
    "1111101110100100",
    "1111101000010101",
    "1111100001100100",
    "1111011010000010",
    "1111010001101011",
    "1111001000100010",
    "1110111110111011",
    "1110110101100100",
    "1110101101001010",
    "1110100110100100",
    "1110100010010010",
    "1110100000101011",
    "1110100001110100",
    "1110100110000000",
    "1110101101100001",
    "1110111000110010",
    "1111000111110010",
    "1111011001100111",
    "1111101100000110",
    "1111111100010010",
    "1111111000110110",
    "1111110101100001",
    "1111111010010010",
    "1111111001110101",
    "1111101001001000",
    "1111010110000011",
    "1111000010100111",
    "1110110000010010",
    "1110011111110110",
    "1110010001111101",
    "1110000111001110",
    "1110000000010101",
    "1101111101110111",
    "1101111111110110",
    "1110000101111011",
    "1110001111010001",
    "1110011011000110",
    "1110101000111001",
    "1110111000011000",
    "1111001001011101",
    "1111011011101111",
    "1111101110010100",
    "1111111111110011",
    "1111110001011100",
    "1111100110110011",
    "1111100000111101",
    "1111011111101100",
    "1111100010010000",
    "1111100111011100",
    "1111101110000100",
    "1111110101001101",
    "1111111100000110",
    "1111111101101111",
    "1111111000111000",
    "1111110101101001",
    "1111110100001111",
    "1111110100101000",
    "1111110110011100",
    "1111111001000101",
    "1111111011111011",
    "1111111110010011",
    "1111111111101110",
    "1111111111111011",
    "1111111110101000",
    "1111111011100001",
    "1111110110010001",
    "1111101110011111",
    "1111100100000110",
    "1111010111011101",
    "1111001001011011",
    "1110111011010011",
    "1110101110011111",
    "1110100100010000",
    "1110011101011001",
    "1110011010010100",
    "1110011011000001",
    "1110011111010110",
    "1110100111010101",
    "1110110011010000",
    "1111000011100010",
    "1111011000011000",
    "1111110001000011",
    "1111110100011010",
    "1111011011001001",
    "1111000110010110",
    "1110111000100101",
    "1110110010110100",
    "1110110100011000",
    "1110111011001111",
    "1111000100111100",
    "1111001111011110",
    "1111011001100011",
    "1111100010101011",
    "1111101010011101",
    "1111110000010100",
    "1111110011010111",
    "1111110010101111",
    "1111101110001100",
    "1111100110011000",
    "1111011100111111",
    "1111010100010101",
    "1111001110100100",
    "1111001101001111",
    "1111010000110011",
    "1111011000101111",
    "1111100100000001",
    "1111110001011111",
    "1111111111111100",
    "1111110001100010",
    "1111100100100101",
    "1111011010100011",
    "1111010100101111",
    "1111010011111110",
    "1111011000011011",
    "1111100001010111",
    "1111101101010111",
    "1111111010101100",
    "1111111000010000",
    "1111101100110001",
    "1111100011011000",
    "1111011100000111",
    "1111010110100010",
    "1111010010000000",
    "1111001101111000",
    "1111001001101101",
    "1111000101010010",
    "1111000000101001",
    "1110111100000001",
    "1110110111110100",
    "1110110100100010",
    "1110110010101001",
    "1110110010011010",
    "1110110011111011",
    "1110110111000001",
    "1110111011100000",
    "1111000001010100",
    "1111001000101100",
    "1111010010010100",
    "1111011111000000",
    "1111101111010101",
    "1111111101000111",
    "1111101000000101",
    "1111010011111100",
    "1111000011010011",
    "1110110111110101",
    "1110110001111110",
    "1110110000111000",
    "1110110010110110",
    "1110110110010011",
    "1110111010101101",
    "1111000000100001",
    "1111001000110111",
    "1111010100100000",
    "1111100011001010",
    "1111110010111110",
    "1111111110111000",
    "1111110101100100",
    "1111110011010110",
    "1111111000101111",
    "1111111011100111",
    "1111101100100011",
    "1111011101010110",
    "1111010000110011",
    "1111001000100010",
    "1111000101000000",
    "1111000101101010",
    "1111001001100010",
    "1111001111100011",
    "1111010110111110",
    "1111011111011001",
    "1111101000100011",
    "1111110010001000",
    "1111111011100101",
    "1111111011111011",
    "1111110101011100",
    "1111110001111011",
    "1111110010000100",
    "1111110110001000",
    "1111111101101110",
    "1111111000001000",
    "1111101100110111",
    "1111100001111110",
    "1111011000110000",
    "1111010010000110",
    "1111001110011100",
    "1111001101110101",
    "1111010000001101",
    "1111010101100100",
    "1111011110000010",
    "1111101001110011",
    "1111111000110111",
    "1111110101001001",
    "1111100001001100",
    "1111001100100011",
    "1110111000110111",
    "1110100111110101",
    "1110011010111101",
    "1110010011001011",
    "1110010000111000",
    "1110010011110001",
    "1110011011000100",
    "1110100101101010",
    "1110110010010111",
    "1111000000001000",
    "1111001110000100",
    "1111011011011101",
    "1111100111101101",
    "1111110010001111",
    "1111111010011110",
    "1111111111111000",
    "1111111101110011",
    "1111111110101001",
    "1111111101101100",
    "1111111000000000",
    "1111110001010011",
    "1111101010110010",
    "1111100101110110",
    "1111100011110011",
    "1111100101110010",
    "1111101100011000",
    "1111110111010001",
    "1111111010110100",
    "1111101100000001",
    "1111011110101001",
    "1111010100101111",
    "1111001111011111",
    "1111001111000100",
    "1111010010100001",
    "1111011000010110",
    "1111011111000111",
    "1111100101110001",
    "1111101100011111",
    "1111110100100110",
    "1111111111111001",
    "1111110000011011",
    "1111011100111101",
    "1111000111111001",
    "1110110100110111",
    "1110100111100111",
    "1110100010101100",
    "1110100110100000",
    "1110110001001000",
    "1110111111000010",
    "1111001100010100",
    "1111010101111100",
    "1111011010011000",
    "1111011001101101",
    "1111010101001101",
    "1111001110101110",
    "1111000111110111",
    "1111000001100110",
    "1110111100010110",
    "1110111000000100",
    "1110110100100101",
    "1110110001101011",
    "1110101111000101",
    "1110101100011110",
    "1110101001011110",
    "1110100101110010",
    "1110100001010010",
    "1110011100000010",
    "1110010110010011",
    "1110010000100100",
    "1110001011011001",
    "1110000111011011",
    "1110000101010010",
    "1110000101011000",
    "1110001000000011",
    "1110001101100011",
    "1110010110001011",
    "1110100010010100",
    "1110110010010100",
    "1111000110001110",
    "1111011101010111",
    "1111110110001110",
    "1111110001100111",
    "1111011100101101",
    "1111001100111100",
    "1111000010111101",
    "1110111110000111",
    "1110111100110010",
    "1110111100111111",
    "1110111101010100",
    "1110111101011110",
    "1110111110001001",
    "1111000000011100",
    "1111000101010010",
    "1111001100011110",
    "1111010100111001",
    "1111011100100101",
    "1111100001100110",
    "1111100010101110",
    "1111011111111000",
    "1111011010001100",
    "1111010011110001",
    "1111001110111010",
    "1111001101101000",
    "1111010001011001",
    "1111011010110010",
    "1111101001011110",
    "1111111100000111",
    "1111101111010010",
    "1111011011001111",
    "1111001001111010",
    "1110111100101110",
    "1110110100010000",
    "1110110000000111",
    "1110101111011100",
    "1110110001011010",
    "1110110101100101",
    "1110111011111100",
    "1111000100101111",
    "1111010000000010",
    "1111011101011011",
    "1111101011111001",
    "1111111010000111",
    "1111111001010100",
    "1111101111100100",
    "1111101001001101",
    "1111100110001101",
    "1111100110000110",
    "1111101000001001",
    "1111101011100110",
    "1111101111101010",
    "1111110011011110",
    "1111110110001011",
    "1111110110110111",
    "1111110100111010",
    "1111101111111111",
    "1111101000010101",
    "1111011110100110",
    "1111010011110011",
    "1111001001000100",
    "1110111111011100",
    "1110110111101000",
    "1110110010000010",
    "1110101110101110",
    "1110101101101101",
    "1110101110111000",
    "1110110010001011",
    "1110110111100111",
    "1110111111001010",
    "1111001000110010",
    "1111010100010101",
    "1111100001010101",
    "1111101111000100",
    "1111111100100000",
    "1111110111100110",
    "1111101110100000",
    "1111101001000111",
    "1111100111110011",
    "1111101010010011",
    "1111101111111011",
    "1111110111101100",
    "1111111111001001",
    "1111110101001111",
    "1111101010110110",
    "1111100000001100",
    "1111010101111011",
    "1111001101001100",
    "1111000111101010",
    "1111000111001101",
    "1111001101001001",
    "1111011001110101",
    "1111101100001111",
    "1111111110000101",
    "1111101000011101",
    "1111010110000110",
    "1111001001011011",
    "1111000011100100",
    "1111000100010000",
    "1111001010001100",
    "1111010011011100",
    "1111011110000100",
    "1111101000010001",
    "1111110000101100",
    "1111110110001111",
    "1111111000001110",
    "1111110110011110",
    "1111110001011010",
    "1111101010001000",
    "1111100010000101",
    "1111011010110101",
    "1111010101100000",
    "1111010010101110",
    "1111010010011100",
    "1111010100000011",
    "1111010110111001",
    "1111011010011001",
    "1111011110011001",
    "1111100010111110",
    "1111101000011000",
    "1111101110110100",
    "1111110110001101",
    "1111111110001001",
    "1111111010000101",
    "1111110011010110",
    "1111101110010101",
    "1111101011010111",
    "1111101010010110",
    "1111101010101111",
    "1111101011110000",
    "1111101100100000",
    "1111101100001010",
    "1111101010000011",
    "1111100101110010",
    "1111011111010111",
    "1111010111000100",
    "1111001101100001",
    "1111000011100110",
    "1110111010010001",
    "1110110010011101",
    "1110101101000000",
    "1110101010100000",
    "1110101011011000",
    "1110101111111111",
    "1110111000011101",
    "1111000100100010",
    "1111010011001010",
    "1111100010100010",
    "1111110000011010",
    "1111111010100000",
    "1111111111001110",
    "1111111110000111",
    "1111110111110011",
    "1111101101110101",
    "1111100010000000",
    "1111010101111110",
    "1111001010110111",
    "1111000001011110",
    "1110111010010110",
    "1110110110000001",
    "1110110100111011",
    "1110110111010001",
    "1110111100111010",
    "1111000101001000",
    "1111001110110000",
    "1111011000011110",
    "1111100001000111",
    "1111100111111011",
    "1111101100100111",
    "1111101111010000",
    "1111101111111111",
    "1111101110110100",
    "1111101011101111",
    "1111100110101010",
    "1111011111110011",
    "1111010111100111",
    "1111001110111000",
    "1111000110100111",
    "1110111111110101",
    "1110111011001111",
    "1110111001010101",
    "1110111010001100",
    "1110111101100000",
    "1111000010101001",
    "1111001000101111",
    "1111001110110000",
    "1111010011101001",
    "1111010110101000",
    "1111010111011000",
    "1111010110000000",
    "1111010011001101",
    "1111001111111010",
    "1111001101000101",
    "1111001011011101",
    "1111001011010110",
    "1111001100110101",
    "1111001111101011",
    "1111010011101001",
    "1111011000011011",
    "1111011101110000",
    "1111100011010111",
    "1111101000111001",
    "1111101110001000",
    "1111110010110101",
    "1111110110111110",
    "1111111010101111",
    "1111111110011001",
    "1111111101110000",
    "1111111001101001",
    "1111110101011010",
    "1111110001010111",
    "1111101110000001",
    "1111101011111000",
    "1111101011010011",
    "1111101100100000",
    "1111101111100010",
    "1111110100011001",
    "1111111011001001",
    "1111111100000111",
    "1111110001100111",
    "1111100101110110",
    "1111011010000100",
    "1111001111110110",
    "1111001000110111",
    "1111000110001101",
    "1111001000000100",
    "1111001101100011",
    "1111010100111011",
    "1111011100001010",
    "1111100001100110",
    "1111100100001110",
    "1111100011111011",
    "1111100001001101",
    "1111011101000100",
    "1111011000100010",
    "1111010100100111",
    "1111010010000011",
    "1111010001011010",
    "1111010011000101",
    "1111010111001001",
    "1111011101100110",
    "1111100110000011",
    "1111110000000011",
    "1111111010110100",
    "1111111010011111",
    "1111110000111000",
    "1111101001001100",
    "1111100100001011",
    "1111100010001010",
    "1111100011000000",
    "1111100110001000",
    "1111101010100010",
    "1111101111000011",
    "1111110010100111",
    "1111110100011111",
    "1111110100001111",
    "1111110001111001",
    "1111101101101011",
    "1111100111111111",
    "1111100001011010",
    "1111011010101000",
    "1111010100011000",
    "1111001111011001",
    "1111001100001001",
    "1111001010111100",
    "1111001011110111",
    "1111001110101101",
    "1111010011001011",
    "1111011000111001",
    "1111011111010110",
    "1111100110000001",
    "1111101100001111",
    "1111110001001111",
    "1111110100001101",
    "1111110100011011",
    "1111110001010011",
    "1111101010011101",
    "1111011111111000",
    "1111010010000101",
    "1111000010001101",
    "1110110010000010",
    "1110100011101001",
    "1110011000111010",
    "1110010011010000",
    "1110010011010111",
    "1110011000111111",
    "1110100011011101",
    "1110110001110001",
    "1111000010111000",
    "1111010101101001",
    "1111101000110010",
    "1111111010101110",
    "1111110110001100",
    "1111101011011100",
    "1111100101101100",
    "1111100100110001",
    "1111100111101000",
    "1111101100101001",
    "1111110010001101",
    "1111110111001101",
    "1111111011010000",
    "1111111110100111",
    "1111111110001010",
    "1111111010100111",
    "1111110110100011",
    "1111110010000110",
    "1111101101100110",
    "1111101001011110",
    "1111100101110111",
    "1111100010110100",
    "1111100000000000",
    "1111011101000000",
    "1111011001011101",
    "1111010101000000",
    "1111001111011111",
    "1111001001000110",
    "1111000010001011",
    "1110111011011011",
    "1110110101101100",
    "1110110001110001",
    "1110110000010001",
    "1110110001010100",
    "1110110100101111",
    "1110111001111001",
    "1110111111111101",
    "1111000110010010",
    "1111001100010110",
    "1111010010000010",
    "1111010111011000",
    "1111011100100011",
    "1111100001101001",
    "1111100110101101",
    "1111101011100111",
    "1111110000010101",
    "1111110100110100",
    "1111111001000100",
    "1111111101000011",
    "1111111111010101",
    "1111111100011000",
    "1111111010011010",
    "1111111001110110",
    "1111111011000110",
    "1111111110101001",
    "1111111011000001",
    "1111110001110101",
    "1111100110001000",
    "1111011000110111",
    "1111001011100101",
    "1111000000000010",
    "1110110111101000",
    "1110110011010000",
    "1110110010111001",
    "1110110101111001",
    "1110111011010001",
    "1111000001110110",
    "1111001000100101",
    "1111001110011110",
    "1111010010100010",
    "1111010011111001",
    "1111010001111110",
    "1111001100110000",
    "1111000100111100",
    "1110111011111100",
    "1110110011100010",
    "1110101101010111",
    "1110101010100011",
    "1110101011010110",
    "1110101111010010",
    "1110110101011010",
    "1110111100100011",
    "1111000011110011",
    "1111001010011110",
    "1111010000001100",
    "1111010100110001",
    "1111011000001110",
    "1111011010101101",
    "1111011100100001",
    "1111011101111011",
    "1111011111010100",
    "1111100000111001",
    "1111100010101110",
    "1111100100100000",
    "1111100101101111",
    "1111100101110001",
    "1111100011111001",
    "1111011111110001",
    "1111011001011101",
    "1111010001100111",
    "1111001001001100",
    "1111000001011001",
    "1110111011001111",
    "1110110111100000",
    "1110110110101000",
    "1110111000101111",
    "1110111101101110",
    "1111000101011011",
    "1111001111110000",
    "1111011100100110",
    "1111101100001101",
    "1111111110101011",
    "1111101100001100",
    "1111010101011010",
    "1110111110101011",
    "1110101010000001",
    "1110011001011001",
    "1110001110000111",
    "1110001000011000",
    "1110000111011101",
    "1110001001111001",
    "1110001110010001",
    "1110010011110001",
    "1110011010100110",
    "1110100011111011",
    "1110110001000101",
    "1111000010110001",
    "1111011000001100",
    "1111101111000011",
    "1111111100000011",
    "1111101100101110",
    "1111100101010101",
    "1111100110011011",
    "1111101110100101",
    "1111111010111111",
    "1111110111100010",
    "1111101011110001",
    "1111100011011111",
    "1111011111010010",
    "1111011110111000",
    "1111100001011010",
    "1111100101111001",
    "1111101011011111",
    "1111110001011101",
    "1111110111001010",
    "1111111100000001",
    "1111111111100101",
    "1111111110010101",
    "1111111101110101",
    "1111111110101010",
    "1111111111010100",
    "1111111100010101",
    "1111111000011000",
    "1111110011011101",
    "1111101101100110",
    "1111100110111011",
    "1111011111110000",
    "1111011000100010",
    "1111010010000000",
    "1111001100111101",
    "1111001010001111",
    "1111001010101000",
    "1111001110011100",
    "1111010101100010",
    "1111011111001101",
    "1111101010010111",
    "1111110101101101",
    "1111111111111001",
    "1111110111010110",
    "1111110001000101",
    "1111101101001001",
    "1111101011010101",
    "1111101011011001",
    "1111101101000111",
    "1111110000011101",
    "1111110101011011",
    "1111111011111011",
    "1111111100001110",
    "1111110011011101",
    "1111101010001011",
    "1111100000110110",
    "1111010111111110",
    "1111010000000111",
    "1111001001110100",
    "1111000101101010",
    "1111000100010111",
    "1111000110010000",
    "1111001011010110",
    "1111010010111110",
    "1111011100000010",
    "1111100101000000",
    "1111101100011111",
    "1111110001100000",
    "1111110011101100",
    "1111110011001000",
    "1111110000001010",
    "1111101011000100",
    "1111100011101100",
    "1111011001101101",
    "1111001101000111",
    "1110111110111010",
    "1110110001000111",
    "1110100110011010",
    "1110100001100010",
    "1110100100100000",
    "1110110000000111",
    "1111000011100100",
    "1111011100100001",
    "1111110111011000",
    "1111101111110011",
    "1111011100101110",
    "1111010001110011",
    "1111001111110110",
    "1111010110000110",
    "1111100010011100",
    "1111110010011011",
    "1111111100000011",
    "1111101010001100",
    "1111011000010000",
    "1111000110000011",
    "1110110011101010",
    "1110100001110100",
    "1110010001101100",
    "1110000100110011",
    "1101111100010111",
    "1101111000111110",
    "1101111010001100",
    "1101111110111101",
    "1110000101111100",
    "1110001110010010",
    "1110010111100101",
    "1110100001111101",
    "1110101101101011",
    "1110111010110111",
    "1111001001010011",
    "1111011000010101",
    "1111100110111011",
    "1111110100000000",
    "1111111110101000",
    "1111111001101110",
    "1111110101001001",
    "1111110011001011",
    "1111110010111111",
    "1111110011100110",
    "1111110100001001",
    "1111110100000010",
    "1111110011001001",
    "1111110001110001",
    "1111110000011110",
    "1111110000000010",
    "1111110001010100",
    "1111110100111001",
    "1111111011000001",
    "1111111100100101",
    "1111110010110001",
    "1111101000100101",
    "1111011111000111",
    "1111010111010001",
    "1111010001100010",
    "1111001101110101",
    "1111001011100000",
    "1111001001101101",
    "1111000111011101",
    "1111000100001011",
    "1110111111100100",
    "1110111001111101",
    "1110110100000011",
    "1110101110110101",
    "1110101011011001",
    "1110101010101010",
    "1110101101001010",
    "1110110011000001",
    "1110111100001001",
    "1111001000001110",
    "1111010110111001",
    "1111100111101110",
    "1111111010001100",
    "1111110010100101",
    "1111011111111111",
    "1111001111011110",
    "1111000010011010",
    "1110111001100111",
    "1110110101000001",
    "1110110011110110",
    "1110110100110111",
    "1110110110110100",
    "1110111000110111",
    "1110111010110111",
    "1110111101000111",
    "1111000000001100",
    "1111000100011000",
    "1111001001101010",
    "1111001111011100",
    "1111010100110001",
    "1111011000101111",
    "1111011010101000",
    "1111011010001110",
    "1111010111110010",
    "1111010100000001",
    "1111001111110011",
    "1111001100000001",
    "1111001001010101",
    "1111001000001000",
    "1111001000100011",
    "1111001010011101",
    "1111001101011110",
    "1111010001001111",
    "1111010101010101",
    "1111011001011101",
    "1111011101010010",
    "1111100000100100",
    "1111100010111110",
    "1111100100001011",
    "1111100011110011",
    "1111100001100110",
    "1111011101011100",
    "1111010111011111",
    "1111010000001010",
    "1111001000001000",
    "1111000000000111",
    "1110111000110100",
    "1110110010101100",
    "1110101101111111",
    "1110101010110100",
    "1110101001001011",
    "1110101001001011",
    "1110101010111100",
    "1110101110100100",
    "1110110100010101",
    "1110111100100110",
    "1111001000010101",
    "1111011000100000",
    "1111101101101100",
    "1111111000101011",
    "1111011100111100",
    "1111000010101110",
    "1110101110000000",
    "1110100001111110",
    "1110011111101110",
    "1110100110000000",
    "1110110001110001",
    "1110111111010100",
    "1111001011100001",
    "1111010100100010",
    "1111011001111001",
    "1111011100000101",
    "1111011100000010",
    "1111011010011001",
    "1111010111101010",
    "1111010100000101",
    "1111010000000000",
    "1111001100001001",
    "1111001001011101",
    "1111001000111100",
    "1111001011011011",
    "1111010001010100",
    "1111011010100011",
    "1111100110101101",
    "1111110100111001",
    "1111111100000101",
    "1111101101110101",
    "1111100001111001",
    "1111011001101000",
    "1111010101100111",
    "1111010101101001",
    "1111011000110000",
    "1111011101101001",
    "1111100011000101",
    "1111101000010001",
    "1111101101000001",
    "1111110001100110",
    "1111110110011011",
    "1111111011101111",
    "1111111110100110",
    "1111111001001001",
    "1111110100101010",
    "1111110001110111",
    "1111110001000110",
    "1111110010010011",
    "1111110100111111",
    "1111111000011001",
    "1111111011101010",
    "1111111110000001",
    "1111111110110110",
    "1111111101110011",
    "1111111010111010",
    "1111110110100111",
    "1111110001101000",
    "1111101100111000",
    "1111101001010000",
    "1111100111011100",
    "1111100111110100",
    "1111101010011000",
    "1111101110110110",
    "1111110100101010",
    "1111111011000011",
    "1111111111000000",
    "1111111010101011",
    "1111111001000110",
    "1111111011000110",
    "1111111110111111",
    "1111110101101100",
    "1111101010001010",
    "1111011110000101",
    "1111010011001010",
    "1111001010100110",
    "1111000101001000",
    "1111000010100111",
    "1111000010100110",
    "1111000100010010",
    "1111000111001000",
    "1111001010101111",
    "1111001111001000",
    "1111010100100100",
    "1111011011010011",
    "1111100011100100",
    "1111101101011011",
    "1111111000100000",
    "1111111011110010",
    "1111110000011000",
    "1111100110000100",
    "1111011101100001",
    "1111010111000011",
    "1111010010011100",
    "1111001111000100",
    "1111001011111101",
    "1111001000000110",
    "1111000010101001",
    "1110111011010110",
    "1110110010100100",
    "1110101001001001",
    "1110100000001100",
    "1110011000101100",
    "1110010011001111",
    "1110010000000010",
    "1110001110111010",
    "1110001111100110",
    "1110010001111110",
    "1110010110000001",
    "1110011011111000",
    "1110100011101110",
    "1110101101100000",
    "1110111000111100",
    "1111000101100000",
    "1111010010100111",
    "1111011111100110",
    "1111101011111110",
    "1111110111010010",
    "1111111110110011",
    "1111110110110111",
    "1111110001001111",
    "1111101110010101",
    "1111101110010101",
    "1111110001001011",
    "1111110110101000",
    "1111111110011000",
    "1111110111111101",
    "1111101100111100",
    "1111100001010100",
    "1111010110001011",
    "1111001100111100",
    "1111000111001001",
    "1111000110001001",
    "1111001010110010",
    "1111010100111110",
    "1111100011100100",
    "1111110100100000",
    "1111111010101101",
    "1111101100101111",
    "1111100011011000",
    "1111011111100011",
    "1111100001000010",
    "1111100110111010",
    "1111101111110100",
    "1111111010011001",
    "1111111010011010",
    "1111101111110000",
    "1111100110101000",
    "1111100000010001",
    "1111011101110101",
    "1111100000001000",
    "1111100111010000",
    "1111110010001110",
    "1111111111001011",
    "1111110100001110",
    "1111101010011010",
    "1111100101001000",
    "1111100101010011",
    "1111101011000011",
    "1111110101111111",
    "1111111010101010",
    "1111101000001110",
    "1111010100010111",
    "1111000001000011",
    "1110110000011001",
    "1110100011111011",
    "1110011100010111",
    "1110011001100011",
    "1110011010011011",
    "1110011101100001",
    "1110100001100110",
    "1110100101111001",
    "1110101010001110",
    "1110101110110110",
    "1110110100000101",
    "1110111010000111",
    "1111000000110110",
    "1111000111111111",
    "1111001111001010",
    "1111010110000100",
    "1111011100101101",
    "1111100011010111",
    "1111101010100001",
    "1111110010111000",
    "1111111101000111",
    "1111110110010101",
    "1111100111101001",
    "1111010111011101",
    "1111000111000011",
    "1110110111110001",
    "1110101010111000",
    "1110100001001101",
    "1110011010111111",
    "1110011000001001",
    "1110011000101000",
    "1110011100110010",
    "1110100101011000",
    "1110110011010000",
    "1111000110110010",
    "1111011111000000",
    "1111111001100010",
    "1111101101001001",
    "1111011000110010",
    "1111001100000101",
    "1111000111111111",
    "1111001011011110",
    "1111010100001000",
    "1111011111000100",
    "1111101001110011",
    "1111110010110111",
    "1111111001101001",
    "1111111101111100",
    "1111111111110001",
    "1111111110111110",
    "1111111011011110",
    "1111110101011101",
    "1111101101100100",
    "1111100100110100",
    "1111011100011011",
    "1111010101011000",
    "1111010000001101",
    "1111001101000000",
    "1111001011100101",
    "1111001011110010",
    "1111001101110011",
    "1111010001111110",
    "1111011000110010",
    "1111100010010010",
    "1111101110001100",
    "1111111011100110",
    "1111110110110000",
    "1111101010011111",
    "1111100001001000",
    "1111011011111111",
    "1111011011110111",
    "1111100000111001",
    "1111101010100111",
    "1111110111110101",
    "1111111001000011",
    "1111101001111010",
    "1111011100010111",
    "1111010001110011",
    "1111001011000010",
    "1111001000010001",
    "1111001001010011",
    "1111001101011110",
    "1111010100000000",
    "1111011100000101",
    "1111100100111110",
    "1111101110000100",
    "1111110110110011",
    "1111111110110011",
    "1111111010000100",
    "1111110011110111",
    "1111101110010101",
    "1111101001001011",
    "1111100100001010",
    "1111011111010001",
    "1111011010110000",
    "1111010111001000",
    "1111010100111011",
    "1111010100011000",
    "1111010101011010",
    "1111010111010110",
    "1111011001010011",
    "1111011010001100",
    "1111011001001011",
    "1111010101100111",
    "1111001111010110",
    "1111000110011010",
    "1110111011010001",
    "1110101110111010",
    "1110100010110110",
    "1110011001000100",
    "1110010011100110",
    "1110010100000101",
    "1110011011010100",
    "1110101000111111",
    "1110111011011001",
    "1111001111110001",
    "1111100010110110",
    "1111110001101010",
    "1111111010000100",
    "1111111011010000",
    "1111110101101100",
    "1111101010111001",
    "1111011100111000",
    "1111001101101101",
    "1110111111001010",
    "1110110010100110",
    "1110101000111010",
    "1110100010100010",
    "1110011111011110",
    "1110011111001111",
    "1110100001000101",
    "1110100100001000",
    "1110100111100000",
    "1110101010101010",
    "1110101101010100",
    "1110101111100011",
    "1110110001101100",
    "1110110100010010",
    "1110110111110101",
    "1110111100110011",
    "1111000011011101",
    "1111001100000010",
    "1111010110010101",
    "1111100001111000",
    "1111101101101000",
    "1111111000001100",
    "1111111111110001",
    "1111111011010011",
    "1111111010100000",
    "1111111100110011",
    "1111111110111001",
    "1111111001110010",
    "1111110100100011",
    "1111101111001000",
    "1111101000101111",
    "1111100000011001",
    "1111010101011000",
    "1111000111111110",
    "1110111001010011",
    "1110101011001111",
    "1110011111110101",
    "1110011000101010",
    "1110010110100100",
    "1110011001110000",
    "1110100010000010",
    "1110101111000010",
    "1111000000000000",
    "1111010011100001",
    "1111100111011000",
    "1111111000110101",
    "1111111010101011",
    "1111110100111110",
    "1111110110100101",
    "1111111110101001",
    "1111110100011100",
    "1111100100101001",
    "1111010011101010",
    "1111000011000011",
    "1110110100010010",
    "1110101000111001",
    "1110100010001010",
    "1110100001001000",
    "1110100101111110",
    "1110101111111011",
    "1110111101011100",
    "1111001100100110",
    "1111011011100101",
    "1111101001010000",
    "1111110100111110",
    "1111111110011010",
    "1111111010101100",
    "1111110111000001",
    "1111110111001000",
    "1111111011011110",
    "1111111100001010",
    "1111110000111000",
    "1111100100010000",
    "1111011000001000",
    "1111001110001001",
    "1111000111010110",
    "1111000100010101",
    "1111000101010000",
    "1111001010000111",
    "1111010010111000",
    "1111011111010010",
    "1111101110101100",
    "1111111111111100",
    "1111101110101000",
    "1111011111000111",
    "1111010011010111",
    "1111001100100110",
    "1111001011001111",
    "1111001110101011",
    "1111010101101001",
    "1111011110101000",
    "1111101000001011",
    "1111110001001110",
    "1111111001000101",
    "1111111111011110",
    "1111111011110000",
    "1111111000100111",
    "1111110111000001",
    "1111110110110001",
    "1111110111101011",
    "1111111001100000",
    "1111111100000100",
    "1111111111001111",
    "1111111100111100",
    "1111111000011111",
    "1111110011010010",
    "1111101101010011",
    "1111100110110010",
    "1111100000010111",
    "1111011011000001",
    "1111010111111100",
    "1111011000010110",
    "1111011101000000",
    "1111100110001101",
    "1111110011001000",
    "1111111101111000",
    "1111101111011011",
    "1111100100001000",
    "1111011110001101",
    "1111011110110110",
    "1111100110000011",
    "1111110010110011",
    "1111111100011001",
    "1111101000111110",
    "1111010011110001",
    "1110111101100011",
    "1110100111011000",
    "1110010010111000",
    "1110000010001000",
    "1101110111000011",
    "1101110010110001",
    "1101110101010010",
    "1101111101001110",
    "1110001000010110",
    "1110010100011000",
    "1110011111011010",
    "1110101000100010",
    "1110101111011110",
    "1110110100100111",
    "1110111000011010",
    "1110111011001110",
    "1110111101011001",
    "1110111111000100",
    "1111000000011001",
    "1111000001100001",
    "1111000010011100",
    "1111000010111110",
    "1111000010110001",
    "1111000001001101",
    "1110111101110101",
    "1110111000011011",
    "1110110001001010",
    "1110101000100111",
    "1110011111100110",
    "1110010111000100",
    "1110001111111101",
    "1110001010110111",
    "1110001000000011",
    "1110000111011011",
    "1110001000110100",
    "1110001011111100",
    "1110010000110000",
    "1110010111011011",
    "1110100000010001",
    "1110101011101111",
    "1110111001111100",
    "1111001010100101",
    "1111011100100001",
    "1111101110000101",
    "1111111101011000",
    "1111110111001010",
    "1111110000010110",
    "1111101101111100",
    "1111101110111001",
    "1111110001101100",
    "1111110100111101",
    "1111110111101011",
    "1111111001011110",
    "1111111010001110",
    "1111111001111011",
    "1111111000011001",
    "1111110101010000",
    "1111110000001000",
    "1111101000110101",
    "1111011111101100",
    "1111010101100100",
    "1111001011110010",
    "1111000011110100",
    "1110111110111111",
    "1110111110001001",
    "1111000001100111",
    "1111001001011011",
    "1111010101001110",
    "1111100100100100",
    "1111110110101111",
    "1111110101001100",
    "1111100000110000",
    "1111001101100100",
    "1110111101010110",
    "1110110001010101",
    "1110101010000110",
    "1110100111011000",
    "1110101000010001",
    "1110101011011110",
    "1110101111101011",
    "1110110011111001",
    "1110110111011011",
    "1110111001110101",
    "1110111010110111",
    "1110111010011001",
    "1110111000100010",
    "1110110101100000",
    "1110110001110001",
    "1110101101111011",
    "1110101010100000",
    "1110100111110001",
    "1110100101101110",
    "1110100100010010",
    "1110100011011100",
    "1110100011110110",
    "1110100110110100",
    "1110101110000000",
    "1110111010101111",
    "1111001101000101",
    "1111100011110110",
    "1111111100011110",
    "1111101100001110",
    "1111011001010001",
    "1111001100011011",
    "1111000101111110",
    "1111000100110001",
    "1111000110111110",
    "1111001010101000",
    "1111001110001111",
    "1111010001000000",
    "1111010010110011",
    "1111010011110110",
    "1111010100011111",
    "1111010101000101",
    "1111010110000001",
    "1111010111101101",
    "1111011010100101",
    "1111011110110001",
    "1111100011111011",
    "1111101001000011",
    "1111101100101011",
    "1111101101001110",
    "1111101001010111",
    "1111100000101001",
    "1111010011101001",
    "1111000100001010",
    "1110110100110001",
    "1110101000001100",
    "1110100000101110",
    "1110011111101100",
    "1110100101100010",
    "1110110001111000",
    "1111000011110100",
    "1111011010001001",
    "1111110010111001",
    "1111110100011000",
    "1111011110101011",
    "1111001110100110",
    "1111000101110110",
    "1111000100101010",
    "1111001001101111",
    "1111010010100010",
    "1111011100010011",
    "1111100100101010",
    "1111101010011000",
    "1111101101001101",
    "1111101101110000",
    "1111101101000000",
    "1111101011110111",
    "1111101010111001",
    "1111101010011100",
    "1111101010101010",
    "1111101011100110",
    "1111101101011010",
    "1111110000000010",
    "1111110011010011",
    "1111110110110110",
    "1111111010011010",
    "1111111101111101",
    "1111111110001101",
    "1111111001101011",
    "1111110011111001",
    "1111101100100000",
    "1111100011100100",
    "1111011001011101",
    "1111001110111111",
    "1111000101000011",
    "1110111100100011",
    "1110110110001101",
    "1110110010010101",
    "1110110001000101",
    "1110110010001010",
    "1110110101001101",
    "1110111001110000",
    "1110111111010010",
    "1111000101011000",
    "1111001011100001",
    "1111010001011010",
    "1111010110111011",
    "1111011100001001",
    "1111100001011111",
    "1111100111100000",
    "1111101110101101",
    "1111110111011001",
    "1111111110100100",
    "1111110100000000",
    "1111101010000110",
    "1111100010010101",
    "1111011110001001",
    "1111011110010001",
    "1111100010110100",
    "1111101011001010",
    "1111110110000100",
    "1111111101110111",
    "1111110010001001",
    "1111100111110100",
    "1111011111100110",
    "1111011001110111",
    "1111010110101111",
    "1111010110000011",
    "1111010111011010",
    "1111011010010011",
    "1111011101111111",
    "1111100001101100",
    "1111100100101111",
    "1111100110101111",
    "1111100111100010",
    "1111100111010011",
    "1111100110010101",
    "1111100100111100",
    "1111100011010101",
    "1111100001100100",
    "1111011111110000",
    "1111011110000010",
    "1111011100110011",
    "1111011100100011",
    "1111011101110111",
    "1111100001010010",
    "1111100111001011",
    "1111101111011101",
    "1111111001100010",
    "1111111011101010",
    "1111110001100110",
    "1111101001100111",
    "1111100100110011",
    "1111100011101111",
    "1111100110100100",
    "1111101100111000",
    "1111110110001000",
    "1111111110010100",
    "1111110001001101",
    "1111100011010101",
    "1111010101101010",
    "1111001001010000",
    "1110111111000111",
    "1110110111110111",
    "1110110011101110",
    "1110110010010010",
    "1110110010110011",
    "1110110100010111",
    "1110110110001001",
    "1110110111110101",
    "1110111001011000",
    "1110111011000111",
    "1110111101101000",
    "1111000001011010",
    "1111000111001110",
    "1111001111101100",
    "1111011011010110",
    "1111101010000110",
    "1111111011001000",
    "1111110011010001",
    "1111100011010000",
    "1111010110110010",
    "1111001110111111",
    "1111001011111100",
    "1111001100110000",
    "1111010000000011",
    "1111010100101111",
    "1111011010010100",
    "1111100001000101",
    "1111101001101001",
    "1111110100011100",
    "1111111110101110",
    "1111110001000100",
    "1111100100010010",
    "1111011001111111",
    "1111010011001000",
    "1111001111011111",
    "1111001101111000",
    "1111001100011110",
    "1111001001110010",
    "1111000100111110",
    "1110111110001101",
    "1110110110011000",
    "1110101110101101",
    "1110101000010101",
    "1110100100000110",
    "1110100010011001",
    "1110100011011000",
    "1110100111010011",
    "1110101110011100",
    "1110111001001001",
    "1111000111101000",
    "1111011001101000",
    "1111101110001010",
    "1111111100010011",
    "1111100111101101",
    "1111010101110110",
    "1111000111111111",
    "1110111110100100",
    "1110111001000111",
    "1110110110100111",
    "1110110101101010",
    "1110110101000001",
    "1110110011110100",
    "1110110001101110",
    "1110101111000100",
    "1110101100011100",
    "1110101010101101",
    "1110101010011110",
    "1110101100001010",
    "1110101111110011",
    "1110110101001011",
    "1110111011111100",
    "1111000011101100",
    "1111001100001001",
    "1111010101001011",
    "1111011110110101",
    "1111101001001000",
    "1111110100000011",
    "1111111111010011",
    "1111110101100100",
    "1111101011010110",
    "1111100010111001",
    "1111011101000000",
    "1111011010100010",
    "1111011011111010",
    "1111100001010101",
    "1111101010011010",
    "1111110110000101",
    "1111111101000101",
    "1111110000111001",
    "1111100111000000",
    "1111100000101001",
    "1111011110011100",
    "1111100000011001",
    "1111100101111011",
    "1111101110000000",
    "1111110111011010",
    "1111111111001000",
    "1111110110111100",
    "1111110000111110",
    "1111101101110100",
    "1111101101101000",
    "1111110000001110",
    "1111110101000111",
    "1111111011110001",
    "1111111100011000",
    "1111110100000110",
    "1111101100001010",
    "1111100101100010",
    "1111100001001111",
    "1111100000000000",
    "1111100010010100",
    "1111101000000110",
    "1111110000111110",
    "1111111100010000",
    "1111110110110101",
    "1111101001010111",
    "1111011100011001",
    "1111010000111101",
    "1111001000000100",
    "1111000010011111",
    "1111000000100011",
    "1111000010001111",
    "1111000111001000",
    "1111001110101000",
    "1111011000000100",
    "1111100010110110",
    "1111101110011000",
    "1111111010001111",
    "1111111001111100",
    "1111101110101001",
    "1111100100010010",
    "1111011011010100",
    "1111010100011101",
    "1111010000010001",
    "1111001111010010",
    "1111010001110110",
    "1111010111111001",
    "1111100001000010",
    "1111101100100011",
    "1111111001110001",
    "1111110111110111",
    "1111101000110011",
    "1111011001011011",
    "1111001010011011",
    "1110111100111010",
    "1110110010010000",
    "1110101011101010",
    "1110101001111010",
    "1110101101000010",
    "1110110100010000",
    "1110111110001111",
    "1111001001010011",
    "1111010011110100",
    "1111011100001110",
    "1111100001001111",
    "1111100010000101",
    "1111011110100100",
    "1111010111011101",
    "1111001110001101",
    "1111000100111011",
    "1110111101101000",
    "1110111001111100",
    "1110111010101101",
    "1110111111110011",
    "1111001000101010",
    "1111010100101100",
    "1111100011101010",
    "1111110101110000",
    "1111110100111110",
    "1111011101011011",
    "1111000101100000",
    "1110110000001100",
    "1110100000101110",
    "1110011001110100",
    "1110011100101101",
    "1110101000111100",
    "1110111100010111",
    "1111010011110100",
    "1111101011101100",
    "1111111111000010",
    "1111101110100010",
    "1111100011101100",
    "1111011110010010",
    "1111011101011001",
    "1111011111100100",
    "1111100011100010",
    "1111101000010010",
    "1111101101010110",
    "1111110010100111",
    "1111111000010100",
    "1111111110110011",
    "1111111001100100",
    "1111110000101111",
    "1111100110110000",
    "1111011011110010",
    "1111010000010001",
    "1111000100101100",
    "1110111001110100",
    "1110110000100001",
    "1110101001101010",
    "1110100101110100",
    "1110100101001011",
    "1110100111010110",
    "1110101011100110",
    "1110110001001000",
    "1110110111001101",
    "1110111101100011",
    "1111000100001010",
    "1111001011001110",
    "1111010010111110",
    "1111011011001111",
    "1111100011101010",
    "1111101011100001",
    "1111110010000011",
    "1111110110100101",
    "1111111000101100",
    "1111111000000110",
    "1111110100101100",
    "1111101110100110",
    "1111100110010000",
    "1111011100101011",
    "1111010011010011",
    "1111001011110011",
    "1111000111100111",
    "1111000111100011",
    "1111001011110010",
    "1111010011110001",
    "1111011110011001",
    "1111101010010110",
    "1111110110000000",
    "1111111111101010",
    "1111111010001010",
    "1111111000110000",
    "1111111100100111",
    "1111111010011001",
    "1111101101000111",
    "1111011100101011",
    "1111001010011011",
    "1110110111110100",
    "1110100110010101",
    "1110010111010001",
    "1110001011101011",
    "1110000100001110",
    "1110000001000111",
    "1110000010000000",
    "1110000110010101",
    "1110001101011001",
    "1110010110100101",
    "1110100001101100",
    "1110101110101000",
    "1110111101010110",
    "1111001101100000",
    "1111011110001100",
    "1111101110000000",
    "1111111011010101",
    "1111111011001000",
    "1111110110001110",
    "1111110101110111",
    "1111111001001000",
    "1111111110100111",
    "1111111011010001",
    "1111110110000000",
    "1111110010100011",
    "1111110001010110",
    "1111110010011001",
    "1111110101001011",
    "1111111001000010",
    "1111111101010010",
    "1111111110101011",
    "1111111011010011",
    "1111111000101111",
    "1111110110111110",
    "1111110101111011",
    "1111110101011101",
    "1111110101100000",
    "1111110110001101",
    "1111110111111001",
    "1111111011000011",
    "1111111111110100",
    "1111111000100101",
    "1111101111011110",
    "1111100101010011",
    "1111011011011001",
    "1111010011001101",
    "1111001110000101",
    "1111001100110111",
    "1111001111110110",
    "1111010110111001",
    "1111100001101011",
    "1111110000000010",
    "1111111101110000",
    "1111100111111000",
    "1111001111010111",
    "1110110110011011",
    "1110100000001111",
    "1110001111111111",
    "1110000111111100",
    "1110001000111111",
    "1110010010100010",
    "1110100011000101",
    "1110111001000110",
    "1111010011000011",
    "1111101111001111",
    "1111110100101001",
    "1111011011101111",
    "1111001000111111",
    "1110111110100110",
    "1110111101001010",
    "1111000011011100",
    "1111001110101001",
    "1111011011100110",
    "1111100111110010",
    "1111110001110010",
    "1111111001011100",
    "1111111111010011",
    "1111111100000101",
    "1111111000101101",
    "1111110111000000",
    "1111110111100010",
    "1111111010100011",
    "1111111111100101",
    "1111111010010000",
    "1111110100010010",
    "1111101111011111",
    "1111101100011001",
    "1111101011000111",
    "1111101011010110",
    "1111101100111001",
    "1111101111011101",
    "1111110010111000",
    "1111110110111100",
    "1111111011011001",
    "1111111111111011",
    "1111111011110100",
    "1111111000001101",
    "1111110101011011",
    "1111110011100010",
    "1111110010011010",
    "1111110001111011",
    "1111110010000000",
    "1111110010101011",
    "1111110011111011",
    "1111110101110000",
    "1111111000000100",
    "1111111010110001",
    "1111111101111101",
    "1111111110000001",
    "1111111000110111",
    "1111110010001111",
    "1111101010010001",
    "1111100001100100",
    "1111011001001011",
    "1111010010010101",
    "1111001110001111",
    "1111001101100110",
    "1111010000100001",
    "1111010110100000",
    "1111011110100011",
    "1111100111100001",
    "1111110000010010",
    "1111111000000100",
    "1111111110011011",
    "1111111100011001",
    "1111110111101001",
    "1111110001111100",
    "1111101010000111",
    "1111011111110001",
    "1111010011100110",
    "1111000111001110",
    "1110111100101101",
    "1110110101110010",
    "1110110011010101",
    "1110110100111011",
    "1110111001000100",
    "1110111101110111",
    "1111000001011100",
    "1111000010100100",
    "1111000000100111",
    "1110111011110000",
    "1110110100101001",
    "1110101100010110",
    "1110100011111001",
    "1110011100001111",
    "1110010110000100",
    "1110010010000000",
    "1110010000100100",
    "1110010010010010",
    "1110010111101100",
    "1110100001000000",
    "1110101110001101",
    "1110111110100011",
    "1111010000101001",
    "1111100010100100",
    "1111110010001001",
    "1111111101100101",
    "1111111100001100",
    "1111111011010011",
    "1111111111000010",
    "1111111001101111",
    "1111110000001100",
    "1111100101001000",
    "1111011000111111",
    "1111001100001110",
    "1110111111010001",
    "1110110010110100",
    "1110100111110101",
    "1110011111010100",
    "1110011001111111",
    "1110011000001110",
    "1110011001111111",
    "1110011110110110",
    "1110100110001110",
    "1110101111101100",
    "1110111010111111",
    "1111001000000100",
    "1111010110101101",
    "1111100110010010",
    "1111110101100001",
    "1111111101011001",
    "1111110100011001",
    "1111110000111110",
    "1111110011110011",
    "1111111100110100",
    "1111110100101100",
    "1111100001111101",
    "1111001100100000",
    "1110110110011011",
    "1110100010001010",
    "1110010010000000",
    "1110000111111001",
    "1110000100101110",
    "1110001000011000",
    "1110010001110001",
    "1110011111011110",
    "1110110000000111",
    "1111000010101100",
    "1111010110010010",
    "1111101001101011",
    "1111111011001110",
    "1111110111000001",
    "1111101111000000",
    "1111101101110111",
    "1111110011101000",
    "1111111110110110",
    "1111110010111110",
    "1111100101000001",
    "1111011010001001",
    "1111010100011100",
    "1111010100111011",
    "1111011011100110",
    "1111100111101010",
    "1111110111101001",
    "1111110110010000",
    "1111100011111110",
    "1111010011010000",
    "1111000101011010",
    "1110111011001111",
    "1110110100111100",
    "1110110010001010",
    "1110110010001010",
    "1110110100000110",
    "1110110111001110",
    "1110111010111010",
    "1110111110101110",
    "1111000010010101",
    "1111000101100101",
    "1111001000010000",
    "1111001010001110",
    "1111001011011001",
    "1111001011110111",
    "1111001011111101",
    "1111001100010001",
    "1111001101100011",
    "1111010000100100",
    "1111010110001001",
    "1111011110111111",
    "1111101011011000",
    "1111111010111100",
    "1111110011101100",
    "1111100010101001",
    "1111010100001010",
    "1111001001111100",
    "1111000100110100",
    "1111000100011100",
    "1111000111100011",
    "1111001100101000",
    "1111010010011100",
    "1111011000011011",
    "1111011110101001",
    "1111100101001110",
    "1111101100000000",
    "1111110010001111",
    "1111110110110001",
    "1111111000011101",
    "1111110110100100",
    "1111110001001111",
    "1111101001011111",
    "1111100000110110",
    "1111011000111111",
    "1111010011001011",
    "1111010000000111",
    "1111001111111111",
    "1111010010101011",
    "1111010111110100",
    "1111011111000000",
    "1111100111110001",
    "1111110001100111",
    "1111111100000010",
    "1111111001100001",
    "1111101111110110",
    "1111100111101010",
    "1111100001100110",
    "1111011110000000",
    "1111011101000000",
    "1111011110010001",
    "1111100001000000",
    "1111100100001011",
    "1111100110100100",
    "1111100110111010",
    "1111100100001000",
    "1111011101100110",
    "1111010011010111",
    "1111000110010000",
    "1110110111101010",
    "1110101001001001",
    "1110011100000100",
    "1110010001010100",
    "1110001001001011",
    "1110000011101010",
    "1110000000101001",
    "1110000000000111",
    "1110000010010100",
    "1110000111100111",
    "1110010000010010",
    "1110011100011001",
    "1110101011100001",
    "1110111100111101",
    "1111001111101001",
    "1111100010011101",
    "1111110100010001",
    "1111111100000001",
    "1111101111100011",
    "1111100111000100",
    "1111100010111011",
    "1111100010111101",
    "1111100110010101",
    "1111101011110110",
    "1111110010001001",
    "1111111000001000",
    "1111111101001101",
    "1111111110100100",
    "1111111010110011",
    "1111110110110001",
    "1111110001111110",
    "1111101100011001",
    "1111100110110010",
    "1111100010011111",
    "1111100001001000",
    "1111100100000011",
    "1111101011100011",
    "1111110110101101",
    "1111111100011110",
    "1111110000101011",
    "1111101000010010",
    "1111100100110100",
    "1111100110100111",
    "1111101100111001",
    "1111110110001110",
    "1111111110111101",
    "1111110100000101",
    "1111101010001010",
    "1111100001111101",
    "1111011100000111",
    "1111011001001100",
    "1111011001101000",
    "1111011101010110",
    "1111100011110001",
    "1111101011101010",
    "1111110011010110",
    "1111111001001000",
    "1111111011100110",
    "1111111010000010",
    "1111110100100000",
    "1111101011111010",
    "1111100001101011",
    "1111010111011000",
    "1111001110011100",
    "1111000111110101",
    "1111000011111001",
    "1111000010010111",
    "1111000010100100",
    "1111000011100010",
    "1111000100010111",
    "1111000100010000",
    "1111000010101100",
    "1110111111100001",
    "1110111010111000",
    "1110110101001110",
    "1110101111001000",
    "1110101001010001",
    "1110100100001011",
    "1110100000011100",
    "1110011110010110",
    "1110011110000111",
    "1110011111110110",
    "1110100011100100",
    "1110101001010001",
    "1110110001000111",
    "1110111011010110",
    "1111001000010001",
    "1111011000000001",
    "1111101010001101",
    "1111111101110011",
    "1111101110111001",
    "1111011110001001",
    "1111010010000110",
    "1111001100011001",
    "1111001101110010",
    "1111010101110110",
    "1111100011010111",
    "1111110100010011",
    "1111111001110001",
    "1111101001100010",
    "1111011101011011",
    "1111010111100011",
    "1111011001010001",
    "1111100010110110",
    "1111110011001010",
    "1111111000001110",
    "1111100010101011",
    "1111001111011100",
    "1111000001000011",
    "1110111000101111",
    "1110110110001011",
    "1110110111111111",
    "1110111100011100",
    "1111000010000011",
    "1111001000010001",
    "1111001111010111",
    "1111011000001001",
    "1111100011010101",
    "1111110001000000",
    "1111111111101011",
    "1111110000011111",
    "1111100011011101",
    "1111011010100110",
    "1111010111001101",
    "1111011001100011",
    "1111100001000011",
    "1111101100010100",
    "1111111001100111",
    "1111111000111011",
    "1111101101001111",
    "1111100100110110",
    "1111100000111110",
    "1111100010001101",
    "1111101000011100",
    "1111110010111111",
    "1111111111011000",
    "1111110000010110",
    "1111100001100001",
    "1111010100010000",
    "1111001001100101",
    "1111000010000110",
    "1110111110000101",
    "1110111101011100",
    "1110111111111010",
    "1111000100111110",
    "1111001011111101",
    "1111010100000101",
    "1111011100100110",
    "1111100101000001",
    "1111101101000111",
    "1111110101000001",
    "1111111101001000",
    "1111111001111100",
    "1111101111110001",
    "1111100100000110",
    "1111010111010110",
    "1111001010100011",
    "1110111111001100",
    "1110110110111011",
    "1110110011000110",
    "1110110100100010",
    "1110111011001001",
    "1111000110001001",
    "1111010011111011",
    "1111100010010010",
    "1111101110111001",
    "1111110111110000",
    "1111111011101110",
    "1111111010101100",
    "1111110101101110",
    "1111101110100010",
    "1111100111001100",
    "1111100001010111",
    "1111011110010001",
    "1111011110011001",
    "1111100010000000",
    "1111101000111110",
    "1111110010111110",
    "1111111111010110",
    "1111110010111100",
    "1111100101010101",
    "1111011001011011",
    "1111010000100111",
    "1111001011110000",
    "1111001010111111",
    "1111001101101110",
    "1111010010111110",
    "1111011001110010",
    "1111100001011001",
    "1111101001011111",
    "1111110010000101",
    "1111111011001101",
    "1111111011001001",
    "1111110001010001",
    "1111100111100010",
    "1111011110011110",
    "1111010110100111",
    "1111010000011001",
    "1111001100000001",
    "1111001001100000",
    "1111001000101100",
    "1111001001010001",
    "1111001011000110",
    "1111001110000111",
    "1111010010011101",
    "1111011000100000",
    "1111100000011001",
    "1111101010000011",
    "1111110100111010",
    "1111111111111011",
    "1111110110000110",
    "1111101110010111",
    "1111101001100101",
    "1111100111110111",
    "1111101000111001",
    "1111101100000101",
    "1111110000111011",
    "1111110111010000",
    "1111111111001010",
    "1111110110111010",
    "1111101010110011",
    "1111011100100110",
    "1111001101001110",
    "1110111110001010",
    "1110110001011100",
    "1110101001000010",
    "1110100110011101",
    "1110101010011001",
    "1110110100011101",
    "1111000011000101",
    "1111010011101100",
    "1111100011011000",
    "1111101111100000",
    "1111110110000110",
    "1111110110011101",
    "1111110000111110",
    "1111100110110011",
    "1111011001010011",
    "1111001001100010",
    "1110111000010110",
    "1110100110111011",
    "1110010110110010",
    "1110001001111111",
    "1110000010011001",
    "1110000001010000",
    "1110000110110001",
    "1110010001111110",
    "1110100001001000",
    "1110110010011101",
    "1111000100100111",
    "1111010110111001",
    "1111101001000011",
    "1111111010110000",
    "1111110100110110",
    "1111100111001110",
    "1111011110000010",
    "1111011010110000",
    "1111011110001001",
    "1111101000000000",
    "1111110111001011",
    "1111110110001011",
    "1111100010010010",
    "1111001111001111",
    "1110111110110101",
    "1110110010011001",
    "1110101010110000",
    "1110101000001011",
    "1110101010010011",
    "1110110000010101",
    "1110111001010101",
    "1111000100001110",
    "1111010000001010",
    "1111011100010100",
    "1111101000010001",
    "1111110011101100",
    "1111111110100000",
    "1111110111010010",
    "1111101101111000",
    "1111100101100000",
    "1111011110100011",
    "1111011001011001",
    "1111010110011000",
    "1111010101100000",
    "1111010110011101",
    "1111011000101010",
    "1111011011011001",
    "1111011110000010",
    "1111100000000010",
    "1111100001000111",
    "1111100001000011",
    "1111011111110101",
    "1111011101010110",
    "1111011001110000",
    "1111010101010000",
    "1111010000001111",
    "1111001011011000",
    "1111000111011011",
    "1111000101010000",
    "1111000101011111",
    "1111001000100111",
    "1111001110111011",
    "1111011000111001",
    "1111100110110111",
    "1111111001010011",
    "1111101111111001",
    "1111010110000110",
    "1110111011111000",
    "1110100100101111",
    "1110010100000101",
    "1110001011111100",
    "1110001100101010",
    "1110010100110100",
    "1110100010000011",
    "1110110010000110",
    "1111000011101100",
    "1111010110011010",
    "1111101010011000",
    "1111111111001011",
    "1111101100010111",
    "1111011010011001",
    "1111001101001001",
    "1111000110000000",
    "1111000101001000",
    "1111001001000001",
    "1111001111010110",
    "1111010101011101",
    "1111011001100010",
    "1111011010110000",
    "1111011001010101",
    "1111010110000000",
    "1111010001100100",
    "1111001100101010",
    "1111000111100010",
    "1111000010100001",
    "1110111101110101",
    "1110111001101111",
    "1110110110011111",
    "1110110100010011",
    "1110110011001111",
    "1110110011001101",
    "1110110100001000",
    "1110110110000110",
    "1110111001011000",
    "1110111110010001",
    "1111000101001000",
    "1111001110010001",
    "1111011001110000",
    "1111100111011111",
    "1111110111000111",
    "1111110111111100",
    "1111100110110010",
    "1111010110101100",
    "1111001001000010",
    "1110111111000000",
    "1110111001001100",
    "1110110111011101",
    "1110111000111010",
    "1110111100010001",
    "1111000000010001",
    "1111000100000011",
    "1111000111011011",
    "1111001010111100",
    "1111001111100001",
    "1111010110001110",
    "1111011111100110",
    "1111101011010000",
    "1111110111110011",
    "1111111100110011",
    "1111110100111011",
    "1111110010011000",
    "1111110110001001",
    "1111111111111001",
    "1111110001000010",
    "1111011111010010",
    "1111001101001010",
    "1110111101001001",
    "1110110001001100",
    "1110101010100101",
    "1110101001101111",
    "1110101110001001",
    "1110110110101100",
    "1111000001110110",
    "1111001110000000",
    "1111011001110100",
    "1111100100010010",
    "1111101101000001",
    "1111110100000110",
    "1111111001111011",
    "1111111111000001",
    "1111111100000110",
    "1111110111001000",
    "1111110001110100",
    "1111101100000001",
    "1111100101100111",
    "1111011110100011",
    "1111010110110001",
    "1111001110010111",
    "1111000101100111",
    "1110111100111000",
    "1110110100101001",
    "1110101101100000",
    "1110100111111010",
    "1110100100001101",
    "1110100010011100",
    "1110100010100100",
    "1110100100101010",
    "1110101001000001",
    "1110110000000111",
    "1110111010100010",
    "1111001000100000",
    "1111011001101000",
    "1111101100101100",
    "1111111111110111",
    "1111101110110000",
    "1111100000110011",
    "1111010110111110",
    "1111010001001101",
    "1111001110101000",
    "1111001110001001",
    "1111001110110110",
    "1111010000000111",
    "1111010001110000",
    "1111010011101111",
    "1111010110010000",
    "1111011001100010",
    "1111011101111111",
    "1111100100001010",
    "1111101100110000",
    "1111111000011100",
    "1111111000011110",
    "1111100110101001",
    "1111010011100111",
    "1111000001111000",
    "1110110100001011",
    "1110101100110011",
    "1110101101000101",
    "1110110101000001",
    "1111000011011010",
    "1111010110000000",
    "1111101001111110",
    "1111111100011001",
    "1111110101001101",
    "1111101100101010",
    "1111101010101101",
    "1111101111010010",
    "1111111001100110",
    "1111110111101011",
    "1111100110011011",
    "1111010100110011",
    "1111000101000110",
    "1110111001011000",
    "1110110011000000",
    "1110110010010000",
    "1110110110100000",
    "1110111110001001",
    "1111000111010101",
    "1111010000011001",
    "1111011000000110",
    "1111011101110011",
    "1111100001001100",
    "1111100010010010",
    "1111100001010000",
    "1111011110001111",
    "1111011001010011",
    "1111010010101001",
    "1111001010101010",
    "1111000001110110",
    "1110111000111110",
    "1110110000101110",
    "1110101001101011",
    "1110100100010000",
    "1110100000101011",
    "1110011111000000",
    "1110011111010100",
    "1110100001011111",
    "1110100101010011",
    "1110101010011000",
    "1110110000010111",
    "1110110110111110",
    "1110111110000000",
    "1111000101011111",
    "1111001101100001",
    "1111010110010101",
    "1111100000001010",
    "1111101011001100",
    "1111110111100111",
    "1111111010101100",
    "1111101100001010",
    "1111011101100000",
    "1111001111101001",
    "1111000011101010",
    "1110111010100000",
    "1110110100110011",
    "1110110010110100",
    "1110110100011000",
    "1110111001000010",
    "1111000000011001",
    "1111001010001011",
    "1111010110100111",
    "1111100101111100",
    "1111111000001100",
    "1111110011011110",
    "1111011110111011",
    "1111001100101110",
    "1110111111011010",
    "1110111000101101",
    "1110111000110101",
    "1110111110011001",
    "1111000110111111",
    "1111001111111111",
    "1111010111011011",
    "1111011100100101",
    "1111011111110110",
    "1111100010010000",
    "1111100101000001",
    "1111101000111011",
    "1111101110001011",
    "1111110100100000",
    "1111111011011001",
    "1111111101100101",
    "1111110110101011",
    "1111101111110110",
    "1111101000111011",
    "1111100001110001",
    "1111011010011011",
    "1111010011000011",
    "1111001011111100",
    "1111000101010111",
    "1110111111101001",
    "1110111011000010",
    "1110110111101101",
    "1110110101110110",
    "1110110101101001",
    "1110110111001001",
    "1110111010100011",
    "1110111111111111",
    "1111000111011111",
    "1111010001001010",
    "1111011100110111",
    "1111101010010111",
    "1111111001001000",
    "1111110111100011",
    "1111101000101101",
    "1111011011010100",
    "1111010000011100",
    "1111001000111001",
    "1111000101001000",
    "1111000101010000",
    "1111001001000010",
    "1111001111111101",
    "1111011001011000",
    "1111100100101111",
    "1111110001100111",
    "1111111111100111",
    "1111110001101100",
    "1111100011001011",
    "1111010101101111",
    "1111001010011101",
    "1111000010010000",
    "1110111101101101",
    "1110111101000010",
    "1111000000001010",
    "1111000110111111",
    "1111010001011100",
    "1111011111000100",
    "1111101110110010",
    "1111111110101110",
    "1111110011011101",
    "1111101010001001",
    "1111100110110101",
    "1111101001101111",
    "1111110001101100",
    "1111111100100100",
    "1111111000001010",
    "1111101110111011",
    "1111101001100000",
    "1111101001001011",
    "1111101110011111",
    "1111111001010110",
    "1111110111000111",
    "1111100100110001",
    "1111010001111000",
    "1111000000111011",
    "1110110100000110",
    "1110101100101010",
    "1110101010110010",
    "1110101101110000",
    "1110110100000011",
    "1110111100001010",
    "1111000100110011",
    "1111001101001110",
    "1111010101001001",
    "1111011100101101",
    "1111100100000001",
    "1111101011001011",
    "1111110010000111",
    "1111111000101000",
    "1111111110100010",
    "1111111100010110",
    "1111111000000100",
    "1111110100011111",
    "1111110001011010",
    "1111101110101000",
    "1111101011111001",
    "1111101001000010",
    "1111100110000001",
    "1111100010111110",
    "1111100000010100",
    "1111011110101101",
    "1111011110110101",
    "1111100001010101",
    "1111100110100000",
    "1111101110001011",
    "1111110111011101",
    "1111111110110110",
    "1111110110001100",
    "1111101111101110",
    "1111101100000110",
    "1111101011011101",
    "1111101101011111",
    "1111110001100110",
    "1111110111010000",
    "1111111110001011",
    "1111111001101111",
    "1111110000100010",
    "1111100110010000",
    "1111011011010100",
    "1111010000100011",
    "1111000111000011",
    "1111000000001010",
    "1110111100111111",
    "1110111101111111",
    "1111000010101110",
    "1111001001110111",
    "1111010001011111",
    "1111010111100101",
    "1111011010011110",
    "1111011001000111",
    "1111010011001101",
    "1111001001000110",
    "1110111011110010",
    "1110101100110111",
    "1110011110000101",
    "1110010001010010",
    "1110000111110100",
    "1110000010010101",
    "1110000000101110",
    "1110000010010000",
    "1110000101110111",
    "1110001010110010",
    "1110010000101001",
    "1110010111101101",
    "1110100000010111",
    "1110101010111000",
    "1110110111000001",
    "1111000011110110",
    "1111001111111011",
    "1111011001100111",
    "1111011111011110",
    "1111100000101011",
    "1111011101000100",
    "1111010101010010",
    "1111001010011000",
    "1110111101111010",
    "1110110001100001",
    "1110100110101111",
    "1110011110111010",
    "1110011010111101",
    "1110011011011001",
    "1110100000010101",
    "1110101001101000",
    "1110110110110111",
    "1111000111011010",
    "1111011010010001",
    "1111101110001100",
    "1111111110011001",
    "1111101101001011",
    "1111011111011100",
    "1111010110000000",
    "1111010000111001",
    "1111001111100011",
    "1111010000111000",
    "1111010011110001",
    "1111010111010011",
    "1111011011000110",
    "1111011111001100",
    "1111100100000101",
    "1111101010001101",
    "1111110001111100",
    "1111111011001001",
    "1111111010101110",
    "1111110000110110",
    "1111101000100001",
    "1111100011001000",
    "1111100001110000",
    "1111100100110100",
    "1111101100000000",
    "1111110110001000",
    "1111111110101010",
    "1111110100110100",
    "1111101110110111",
    "1111101110111010",
    "1111110110010001",
    "1111111011000001",
    "1111100110101000",
    "1111001111010100",
    "1110111000101000",
    "1110100110000000",
    "1110011001111100",
    "1110010101100111",
    "1110011000011110",
    "1110100000110110",
    "1110101100010001",
    "1110111000011000",
    "1111000011011101",
    "1111001100101000",
    "1111010100001101",
    "1111011011010001",
    "1111100011000101",
    "1111101100100010",
    "1111110111100101",
    "1111111100100110",
    "1111110001011111",
    "1111101000011100",
    "1111100010001011",
    "1111011110100001",
    "1111011100100000",
    "1111011010110010",
    "1111011000010001",
    "1111010100100100",
    "1111001111111011",
    "1111001011001110",
    "1111000111010101",
    "1111000100110111",
    "1111000011111110",
    "1111000100010111",
    "1111000101011011",
    "1111000110101000",
    "1111000111100101",
    "1111001000000110",
    "1111001000001001",
    "1111000111100111",
    "1111000110011111",
    "1111000100100101",
    "1111000001111001",
    "1110111110011111",
    "1110111010101010",
    "1110110110110010",
    "1110110011100100",
    "1110110001101100",
    "1110110001111000",
    "1110110100110100",
    "1110111011000100",
    "1111000101000001",
    "1111010010101011",
    "1111100011010101",
    "1111110101100000",
    "1111111000111100",
    "1111101010010010",
    "1111100000010100",
    "1111011011110011",
    "1111011100101000",
    "1111100001110000",
    "1111101001111000",
    "1111110011111110",
    "1111111111011111",
    "1111110011110010",
    "1111100110010010",
    "1111011000111100",
    "1111001101100000",
    "1111000110001001",
    "1111000100111011",
    "1111001011000010",
    "1111011000001110",
    "1111101010100110",
    "1111111111000101",
    "1111101101110010",
    "1111011110110110",
    "1111010101101111",
    "1111010010100111",
    "1111010100101001",
    "1111011010011001",
    "1111100010101011",
    "1111101100101010",
    "1111111000001100",
    "1111111010100000",
    "1111101011010111",
    "1111011010101010",
    "1111001001010110",
    "1110111001001011",
    "1110101100001111",
    "1110100100100111",
    "1110100011110011",
    "1110101010001110",
    "1110110111000100",
    "1111001000010110",
    "1111011011010110",
    "1111101101001111",
    "1111111011110001",
    "1111111010010010",
    "1111110101001111",
    "1111110100011001",
    "1111110110110000",
    "1111111011010011",
    "1111111110101001",
    "1111110111100100",
    "1111101111110100",
    "1111100111101111",
    "1111100000000000",
    "1111011001010101",
    "1111010100100000",
    "1111010010001101",
    "1111010010110011",
    "1111010110010000",
    "1111011100011001",
    "1111100100101111",
    "1111101110100110",
    "1111111001001011",
    "1111111100011001",
    "1111110011001001",
    "1111101011111011",
    "1111100111100010",
    "1111100110011110",
    "1111101001000100",
    "1111101111011011",
    "1111111001100110",
    "1111111000100000",
    "1111100111010100",
    "1111010011101010",
    "1110111111000100",
    "1110101011010100",
    "1110011010011101",
    "1110001101111010",
    "1110000110100000",
    "1110000100001011",
    "1110000110001001",
    "1110001011001110",
    "1110010010010100",
    "1110011010101010",
    "1110100011111100",
    "1110101110000101",
    "1110111000101111",
    "1111000011000001",
    "1111001011100101",
    "1111010000100111",
    "1111010000110000",
    "1111001011011011",
    "1111000001010111",
    "1110110100011100",
    "1110100111001000",
    "1110011011111100",
    "1110010100110110",
    "1110010010111110",
    "1110010110110010",
    "1110100000001000",
    "1110101110100100",
    "1111000001010100",
    "1111010111001000",
    "1111101110001001",
    "1111111011111110",
    "1111101001101100",
    "1111011100110010",
    "1111010101111011",
    "1111010100100010",
    "1111010111000110",
    "1111011011101000",
    "1111100000011100",
    "1111100100101001",
    "1111101000000110",
    "1111101011001110",
    "1111101110101000",
    "1111110010110100",
    "1111111000000101",
    "1111111110100011",
    "1111111001110010",
    "1111110001001111",
    "1111101000010010",
    "1111011111101100",
    "1111011000011101",
    "1111010011011111",
    "1111010001011110",
    "1111010010100001",
    "1111010110001101",
    "1111011011101000",
    "1111100001111000",
    "1111101000001110",
    "1111101110011011",
    "1111110100101011",
    "1111111011011011",
    "1111111100111110",
    "1111110100100101",
    "1111101011110011",
    "1111100011100100",
    "1111011100111101",
    "1111011001000110",
    "1111011000111001",
    "1111011101000000",
    "1111100101100100",
    "1111110001110111",
    "1111111111100011",
    "1111110000111010",
    "1111100100100000",
    "1111011100010110",
    "1111011001101000",
    "1111011100011011",
    "1111100011111011",
    "1111101110110100",
    "1111111011110111",
    "1111110101110001",
    "1111100110100101",
    "1111010110101101",
    "1111000110011101",
    "1110110110100100",
    "1110101000010101",
    "1110011101100000",
    "1110010111100111",
    "1110010111011111",
    "1110011100111111",
    "1110100110110110",
    "1110110011010010",
    "1111000000010111",
    "1111001100011011",
    "1111010110100000",
    "1111011110000100",
    "1111100011000110",
    "1111100101110010",
    "1111100110011101",
    "1111100101011000",
    "1111100010111101",
    "1111011111101000",
    "1111011100000101",
    "1111011001001011",
    "1111010111110010",
    "1111011000101111",
    "1111011100100001",
    "1111100011001010",
    "1111101100000100",
    "1111110110011011",
    "1111111110110101",
    "1111110100110100",
    "1111101100010101",
    "1111100101111011",
    "1111100001110100",
    "1111100000000011",
    "1111100000100001",
    "1111100011000001",
    "1111100111011000",
    "1111101101010001",
    "1111110100010101",
    "1111111100000010",
    "1111111100000100",
    "1111110100100001",
    "1111101101101000",
    "1111100111100010",
    "1111100010010111",
    "1111011110001100",
    "1111011011001010",
    "1111011001101000",
    "1111011001110111",
    "1111011100001100",
    "1111100000101011",
    "1111100111000111",
    "1111101110111010",
    "1111110111000111",
    "1111111110101011",
    "1111111011011001",
    "1111110111110111",
    "1111110110111111",
    "1111111000101011",
    "1111111100100010",
    "1111111101101110",
    "1111110110011001",
    "1111101101011000",
    "1111100010010101",
    "1111010101000101",
    "1111000110000110",
    "1110110110101100",
    "1110101000110100",
    "1110011110100100",
    "1110011001100011",
    "1110011010011000",
    "1110100000010100",
    "1110101001100101",
    "1110110011111000",
    "1110111100111111",
    "1111000011010010",
    "1111000101110111",
    "1111000100101001",
    "1111000000000011",
    "1110111001000010",
    "1110110000110101",
    "1110101000110101",
    "1110100010011101",
    "1110011110111111",
    "1110011111001111",
    "1110100011101001",
    "1110101011111010",
    "1110110111010000",
    "1111000100011100",
    "1111010010001000",
    "1111011111000100",
    "1111101010010000",
    "1111110011000110",
    "1111111001100001",
    "1111111101111110",
    "1111111110101001",
    "1111111011011001",
    "1111110111010111",
    "1111110010000110",
    "1111101011101110",
    "1111100100110110",
    "1111011110010111",
    "1111011001010110",
    "1111010110100010",
    "1111010110010011",
    "1111011000101101",
    "1111011101011110",
    "1111100100001011",
    "1111101100011110",
    "1111110110001100",
    "1111111110101001",
    "1111110010000100",
    "1111100100010010",
    "1111010101110100",
    "1111000111101111",
    "1110111011001100",
    "1110110001010010",
    "1110101010110010",
    "1110100111111100",
    "1110101000101000",
    "1110101100100101",
    "1110110011100111",
    "1110111101111000",
    "1111001011101011",
    "1111011101000101",
    "1111110001011110",
    "1111111000111101",
    "1111100100111100",
    "1111010101011010",
    "1111001100100101",
    "1111001011010100",
    "1111010000110000",
    "1111011010101011",
    "1111100110001011",
    "1111110000101000",
    "1111111000010100",
    "1111111100100111",
    "1111111101110001",
    "1111111100100001",
    "1111111001101010",
    "1111110101111000",
    "1111110001101010",
    "1111101101011001",
    "1111101001011111",
    "1111100110011000",
    "1111100100100100",
    "1111100100010010",
    "1111100101101111",
    "1111101000110001",
    "1111101101001101",
    "1111110010101100",
    "1111111000111000",
    "1111111111001101",
    "1111111011000001",
    "1111110110110000",
    "1111110100110100",
    "1111110101111011",
    "1111111010011000",
    "1111111101111111",
    "1111110011111001",
    "1111101000001111",
    "1111011100000001",
    "1111010000000011",
    "1111000100111110",
    "1110111010111100",
    "1110110010000101",
    "1110101010010110",
    "1110100011110100",
    "1110011110101001",
    "1110011011000111",
    "1110011001011011",
    "1110011001101111",
    "1110011100000001",
    "1110100000000111",
    "1110100101110010",
    "1110101100110000",
    "1110110100110001",
    "1110111101101101",
    "1111000111100000",
    "1111010010010000",
    "1111011110000000",
    "1111101010110000",
    "1111111000010011",
    "1111111001110001",
    "1111101100010111",
    "1111100000011100",
    "1111010111000011",
    "1111010000111001",
    "1111001110001100",
    "1111001110011100",
    "1111010000101100",
    "1111010011011101",
    "1111010101001110",
    "1111010100101110",
    "1111010001001100",
    "1111001010101101",
    "1111000010000011",
    "1110111000100101",
    "1110101111110110",
    "1110101001010011",
    "1110100101110110",
    "1110100101110001",
    "1110101000101100",
    "1110101101110111",
    "1110110100011100",
    "1110111011111101",
    "1111000100010000",
    "1111001101011100",
    "1111010111100101",
    "1111100010010111",
    "1111101101000100",
    "1111110110101111",
    "1111111110100001",
    "1111111011111000",
    "1111111000010001",
    "1111110101110111",
    "1111110011111000",
    "1111110001101111",
    "1111101111010111",
    "1111101100111110",
    "1111101011000110",
    "1111101010001000",
    "1111101010010100",
    "1111101011101101",
    "1111101110001111",
    "1111110001111000",
    "1111110110100111",
    "1111111100011000",
    "1111111101001010",
    "1111110110111010",
    "1111110010000001",
    "1111101111110111",
    "1111110001100010",
    "1111110111100000",
    "1111111110100000",
    "1111110001100000",
    "1111100010110110",
    "1111010100000101",
    "1111000110100111",
    "1110111011110000",
    "1110110100100000",
    "1110110001100110",
    "1110110011100001",
    "1110111010100000",
    "1111000110100101",
    "1111010111010011",
    "1111101011100011",
    "1111111110011110",
    "1111101001000010",
    "1111010110010011",
    "1111000111111100",
    "1110111110101101",
    "1110111010011000",
    "1110111010000001",
    "1110111100010001",
    "1110111111110011",
    "1111000011100111",
    "1111000111011000",
    "1111001011011011",
    "1111010000011111",
    "1111010111010011",
    "1111100000000010",
    "1111101010000101",
    "1111110100000011",
    "1111111100001101",
    "1111111110111001",
    "1111111101111010",
    "1111111111011111",
    "1111111010110010",
    "1111110101110001",
    "1111110010010111",
    "1111110010000000",
    "1111110101100010",
    "1111111101000100",
    "1111110111101011",
    "1111101001011001",
    "1111011000111111",
    "1111000111100010",
    "1110110110011010",
    "1110100111000110",
    "1110011010111111",
    "1110010011000110",
    "1110001111110101",
    "1110010000111011",
    "1110010101110001",
    "1110011101100110",
    "1110100111101111",
    "1110110011101100",
    "1111000001000101",
    "1111001111101000",
    "1111011110111011",
    "1111101110011110",
    "1111111101011111",
    "1111110100111010",
    "1111101001110010",
    "1111100001111001",
    "1111011101100110",
    "1111011100111000",
    "1111011111010111",
    "1111100100011000",
    "1111101011010100",
    "1111110011100110",
    "1111111100110100",
    "1111111001001101",
    "1111101110101111",
    "1111100011111100",
    "1111011001010011",
    "1111001111101000",
    "1111000111110111",
    "1111000011000000",
    "1111000001101100",
    "1111000100001000",
    "1111001001110111",
    "1111010001111000",
    "1111011010110100",
    "1111100011001010",
    "1111101001100011",
    "1111101101000101",
    "1111101101010000",
    "1111101001111101",
    "1111100011011000",
    "1111011010000001",
    "1111001110110000",
    "1111000010111110",
    "1110111000100011",
    "1110110001010111",
    "1110101111000111",
    "1110110010110110",
    "1110111101000100",
    "1111001101011110",
    "1111100011000011",
    "1111111011110110",
    "1111101010101111",
    "1111010011101110",
    "1111000001101100",
    "1110110110010011",
    "1110110001111011",
    "1110110011101110",
    "1110111001111111",
    "1111000011000011",
    "1111001101101110",
    "1111011001101111",
    "1111100111001011",
    "1111110110010111",
    "1111111000110010",
    "1111100111000011",
    "1111010101100111",
    "1111000101111110",
    "1110111001010110",
    "1110110000011110",
    "1110101011011011",
    "1110101001111100",
    "1110101011011001",
    "1110101111010100",
    "1110110101000110",
    "1110111100001010",
    "1111000011110110",
    "1111001011100001",
    "1111010010101100",
    "1111011001001001",
    "1111011110110001",
    "1111100011101010",
    "1111100111111001",
    "1111101011011111",
    "1111101110010100",
    "1111110000010000",
    "1111110001000110",
    "1111110000110011",
    "1111101111011111",
    "1111101101100001",
    "1111101011010101",
    "1111101001011110",
    "1111101000010010",
    "1111101000000000",
    "1111101000101101",
    "1111101010011001",
    "1111101101000000",
    "1111110000011111",
    "1111110100101011",
    "1111111001010011",
    "1111111101111010",
    "1111111101111111",
    "1111111011000101",
    "1111111001111100",
    "1111111011001001",
    "1111111111000111",
    "1111111001110110",
    "1111101111111111",
    "1111100011111001",
    "1111010110101101",
    "1111001001111111",
    "1110111111011111",
    "1110111000101101",
    "1110110110100101",
    "1110111001010001",
    "1111000000010100",
    "1111001010110100",
    "1111010111110111",
    "1111100110110110",
    "1111110111101011",
    "1111110101100000",
    "1111100000111110",
    "1111001011101011",
    "1110110111010101",
    "1110100101111110",
    "1110011001100010",
    "1110010011000110",
    "1110010010101111",
    "1110010111101010",
    "1110100000100100",
    "1110101100100001",
    "1110111010111111",
    "1111001011110111",
    "1111011110110001",
    "1111110010111000",
    "1111111001011111",
    "1111101000011111",
    "1111011011111111",
    "1111010100111110",
    "1111010011010000",
    "1111010101011011",
    "1111011001011110",
    "1111011101011011",
    "1111011111110011",
    "1111100000000010",
    "1111011110010001",
    "1111011011000010",
    "1111010110111110",
    "1111010010101001",
    "1111001110011111",
    "1111001010110100",
    "1111000111110111",
    "1111000101110111",
    "1111000101000110",
    "1111000101101110",
    "1111000111110111",
    "1111001011100001",
    "1111010000101001",
    "1111010111001000",
    "1111011110110011",
    "1111100111011000",
    "1111110000100101",
    "1111111010000110",
    "1111111100000011",
    "1111110001101111",
    "1111100110100100",
    "1111011010010011",
    "1111001101001100",
    "1110111111111010",
    "1110110011100100",
    "1110101001101010",
    "1110100011100010",
    "1110100010001011",
    "1110100110000000",
    "1110101110101110",
    "1110111011011001",
    "1111001010011110",
    "1111011001111101",
    "1111100111110001",
    "1111110010000101",
    "1111110111101010",
    "1111110111111100",
    "1111110010111110",
    "1111101001001110",
    "1111011011100001",
    "1111001011000100",
    "1110111001011000",
    "1110101000010001",
    "1110011001101011",
    "1110001111010010",
    "1110001010001011",
    "1110001010100011",
    "1110001111110000",
    "1110011000011000",
    "1110100010101111",
    "1110101101000100",
    "1110110101110111",
    "1110111011111101",
    "1110111110100100",
    "1110111101011100",
    "1110111000111001",
    "1110110001101011",
    "1110101001000100",
    "1110100000101011",
    "1110011001111111",
    "1110010110010000",
    "1110010110000011",
    "1110011001011101",
    "1110100000000000",
    "1110101001000100",
    "1110110011111011",
    "1111000000000011",
    "1111001100111111",
    "1111011010010100",
    "1111100111100101",
    "1111110100001110",
    "1111111111100010",
    "1111110111001000",
    "1111110000011000",
    "1111101100011000",
    "1111101011000000",
    "1111101011110101",
    "1111101110010011",
    "1111110001110110",
    "1111110110000101",
    "1111111010110001",
    "1111111111111001",
    "1111111010011101",
    "1111110100010000",
    "1111101101011101",
    "1111100110000011",
    "1111011101111111",
    "1111010101001110",
    "1111001011101101",
    "1111000001011100",
    "1110110110101111",
    "1110101100001111",
    "1110100010111000",
    "1110011011101011",
    "1110010111100101",
    "1110010111001000",
    "1110011010010110",
    "1110100000111011",
    "1110101010010001",
    "1110110101111001",
    "1111000011011100",
    "1111010010100001",
    "1111100010100001",
    "1111110010011110",
    "1111111111000110",
    "1111110011110110",
    "1111101101000011",
    "1111101011001111",
    "1111101110000011",
    "1111110100011101",
    "1111111101000000",
    "1111111001100010",
    "1111110000010010",
    "1111100111110110",
    "1111100000101011",
    "1111011011000010",
    "1111010111001000",
    "1111010100111100",
    "1111010100010111",
    "1111010100111110",
    "1111010110010011",
    "1111010111111110",
    "1111011001101011",
    "1111011011010011",
    "1111011100110101",
    "1111011110010100",
    "1111011111100100",
    "1111100000010111",
    "1111100000011001",
    "1111011111011111",
    "1111011101110010",
    "1111011011101011",
    "1111011001110111",
    "1111011001001011",
    "1111011010010100",
    "1111011101110101",
    "1111100100000000",
    "1111101100101110",
    "1111110111101010",
    "1111111011110011",
    "1111101110100010",
    "1111100001010111",
    "1111010101000110",
    "1111001010011101",
    "1111000001111000",
    "1110111011101101",
    "1110111000000011",
    "1110110110110010",
    "1110110111110010",
    "1110111010111010",
    "1110111111111111",
    "1111000110111001",
    "1111001111100011",
    "1111011001101011",
    "1111100100111110",
    "1111110000110001",
    "1111111100010101",
    "1111111001001101",
    "1111110000110110",
    "1111101011010000",
    "1111101000111000",
    "1111101001111100",
    "1111101110010100",
    "1111110101101111",
    "1111111111101110",
    "1111110100011001",
    "1111100111110000",
    "1111011011101011",
    "1111010001110110",
    "1111001011110111",
    "1111001010111100",
    "1111001111011110",
    "1111011000110100",
    "1111100101001110",
    "1111110010001111",
    "1111111101001101",
    "1111111100000000",
    "1111111010110000",
    "1111111111011001",
    "1111110110100000",
    "1111100111110110",
    "1111010101101010",
    "1111000001010100",
    "1110101100100110",
    "1110011001101010",
    "1110001010110010",
    "1110000001110000",
    "1101111111011110",
    "1110000011110001",
    "1110001101001110",
    "1110011001110010",
    "1110100111010000",
    "1110110011110100",
    "1110111110001111",
    "1111000101111001",
    "1111001010101011",
    "1111001100110011",
    "1111001100100101",
    "1111001010011110",
    "1111000111001011",
    "1111000011011100",
    "1111000000001010",
    "1110111110000100",
    "1110111101100110",
    "1110111110101011",
    "1111000000111000",
    "1111000011100100",
    "1111000110000110",
    "1111001000000100",
    "1111001001011000",
    "1111001010001001",
    "1111001010101111",
    "1111001011100001",
    "1111001100110010",
    "1111001110100100",
    "1111010000110000",
    "1111010011000011",
    "1111010101010011",
    "1111010111011101",
    "1111011001110000",
    "1111011100101010",
    "1111100000101100",
    "1111100110011110",
    "1111101110010000",
    "1111110111111101",
    "1111111100110111",
    "1111110001000101",
    "1111100101101110",
    "1111011011101011",
    "1111010011101001",
    "1111001101111011",
    "1111001010100101",
    "1111001001011101",
    "1111001010101111",
    "1111001110110000",
    "1111010110001000",
    "1111100001010000",
    "1111110000000000",
    "1111111110100111",
    "1111101100100010",
    "1111011100000101",
    "1111001111011001",
    "1111000111100101",
    "1111000100011111",
    "1111000100110011",
    "1111000110100101",
    "1111000111111110",
    "1111000111110001",
    "1111000101101001",
    "1111000010000010",
    "1110111101101011",
    "1110111001010001",
    "1110110101001011",
    "1110110001010000",
    "1110101101010100",
    "1110101001000010",
    "1110100100010101",
    "1110011111011010",
    "1110011010101111",
    "1110010110111011",
    "1110010100101001",
    "1110010100100100",
    "1110010111001001",
    "1110011100101101",
    "1110100101010111",
    "1110110000110001",
    "1110111110011001",
    "1111001101011100",
    "1111011101000100",
    "1111101100100000",
    "1111111011000110",
    "1111110111101011",
    "1111101100100000",
    "1111100011110100",
    "1111011110000100",
    "1111011011011000",
    "1111011011011110",
    "1111011101101011",
    "1111100000111001",
    "1111100100000101",
    "1111100110010110",
    "1111100111011000",
    "1111100111010100",
    "1111100110110010",
    "1111100110100000",
    "1111100111000100",
    "1111101000101101",
    "1111101011010001",
    "1111101110011000",
    "1111110001100100",
    "1111110100011101",
    "1111110110111001",
    "1111111000111110",
    "1111111011000010",
    "1111111101100101",
    "1111111110110111",
    "1111111010000011",
    "1111110011111100",
    "1111101101000001",
    "1111100110000000",
    "1111011111101110",
    "1111011010111100",
    "1111011000001011",
    "1111010111101000",
    "1111011001010101",
    "1111011101001111",
    "1111100011011111",
    "1111101100001010",
    "1111110111001011",
    "1111111011111010",
    "1111101110001011",
    "1111100001001100",
    "1111010110101101",
    "1111010000011010",
    "1111001111010010",
    "1111010011001101",
    "1111011011000010",
    "1111100100101100",
    "1111101101101101",
    "1111110011101111",
    "1111110101001011",
    "1111110001011110",
    "1111101001001101",
    "1111011101111101",
    "1111010001110001",
    "1111000110110100",
    "1110111110110001",
    "1110111010100101",
    "1110111010010110",
    "1110111101011011",
    "1111000010101011",
    "1111001000110100",
    "1111001110101000",
    "1111010011001011",
    "1111010101111011",
    "1111010110101101",
    "1111010101110010",
    "1111010011101100",
    "1111010001001010",
    "1111001111001010",
    "1111001110101001",
    "1111010000011001",
    "1111010100111110",
    "1111011100100001",
    "1111100110110010",
    "1111110010111101",
    "1111111111111001",
    "1111110011101010",
    "1111101000111110",
    "1111100000110011",
    "1111011011011101",
    "1111011000110000",
    "1111011000001100",
    "1111011001000110",
    "1111011011000001",
    "1111011101110111",
    "1111100001111101",
    "1111101000000010",
    "1111110000111110",
    "1111111101010000",
    "1111110011011000",
    "1111100010010101",
    "1111010001100111",
    "1111000011100110",
    "1110111010001111",
    "1110110110110001",
    "1110111001010101",
    "1111000001011001",
    "1111001101110000",
    "1111011100110101",
    "1111101100101111",
    "1111111011010010",
    "1111111001110000",
    "1111110100010110",
    "1111110101100010",
    "1111111101010101",
    "1111110101010101",
    "1111100100011101",
    "1111010010010101",
    "1111000001001010",
    "1110110010110011",
    "1110101000011110",
    "1110100010111001",
    "1110100010001101",
    "1110100110010110",
    "1110101111000000",
    "1110111011101000",
    "1111001011010110",
    "1111011100111101",
    "1111101110111101",
    "1111111111110011",
    "1111110001111100",
    "1111100111010100",
    "1111100000110011",
    "1111011110011100",
    "1111011111111010",
    "1111100100101111",
    "1111101100011011",
    "1111110110011010",
    "1111111101111110",
    "1111110001110000",
    "1111100110001000",
    "1111011100011110",
    "1111010110001110",
    "1111010100010101",
    "1111010111001101",
    "1111011110011100",
    "1111101001000010",
    "1111110101100010",
    "1111111101100100",
    "1111110001101010",
    "1111100111110000",
    "1111100000011110",
    "1111011100000010",
    "1111011010011000",
    "1111011011001100",
    "1111011110000000",
    "1111100010010100",
    "1111100111101010",
    "1111101101101111",
    "1111110100011010",
    "1111111011101100",
    "1111111100010011",
    "1111110011100110",
    "1111101010010111",
    "1111100001001000",
    "1111011000110010",
    "1111010010011010",
    "1111001111000000",
    "1111001111010001",
    "1111010011011010",
    "1111011011001010",
    "1111100101101010",
    "1111110001100010",
    "1111111101000001",
    "1111111001110010",
    "1111110100101110",
    "1111110101001101",
    "1111111100000010",
    "1111110110110011",
    "1111100100011100",
    "1111001110111000",
    "1110111000111111",
    "1110100101101010",
    "1110010111011101",
    "1110001111110110",
    "1110001111001000",
    "1110010100100000",
    "1110011110100001",
    "1110101011101101",
    "1110111010110101",
    "1111001010111100",
    "1111011011010011",
    "1111101011000111",
    "1111111001011001",
    "1111111010101101",
    "1111110010000001",
    "1111101100101010",
    "1111101010001010",
    "1111101001100010",
    "1111101001100010",
    "1111101001000100",
    "1111100111100001",
    "1111100100110111",
    "1111100001100001",
    "1111011110000101",
    "1111011010111100",
    "1111011000011000",
    "1111010110011010",
    "1111010100111110",
    "1111010100000000",
    "1111010011100010",
    "1111010011101010",
    "1111010100011101",
    "1111010101110100",
    "1111010111100111",
    "1111011001100111",
    "1111011011100000",
    "1111011101001100",
    "1111011110101000",
    "1111011111111011",
    "1111100001010100",
    "1111100010111011",
    "1111100100111001",
    "1111100111001110",
    "1111101001111110",
    "1111101101001111",
    "1111110001001110",
    "1111110110001110",
    "1111111100100111",
    "1111111011011010",
    "1111110001111101",
    "1111100111100010",
    "1111011101001110",
    "1111010100010010",
    "1111001110001100",
    "1111001011111101",
    "1111001110001111",
    "1111010101000101",
    "1111100000000101",
    "1111101110011010",
    "1111111110110010",
    "1111110000011100",
    "1111100001010111",
    "1111010101110001",
    "1111001111000100",
    "1111001101110011",
    "1111010001100111",
    "1111011001100000",
    "1111100100001110",
    "1111110000110001",
    "1111111110100001",
    "1111110010111100",
    "1111100100001011",
    "1111010110001000",
    "1111001010000001",
    "1111000001010101",
    "1110111101000101",
    "1110111101101101",
    "1111000010101110",
    "1111001011001001",
    "1111010101101110",
    "1111100001010101",
    "1111101101001010",
    "1111111000011100",
    "1111111101101001",
    "1111110110010001",
    "1111110010011111",
    "1111110011001001",
    "1111111000011011",
    "1111111110011010",
    "1111110010111110",
    "1111100111001100",
    "1111011101000010",
    "1111010101111110",
    "1111010010101011",
    "1111010011000110",
    "1111010110110001",
    "1111011100110010",
    "1111100100010010",
    "1111101100011001",
    "1111110100010110",
    "1111111011011001",
    "1111111111000110",
    "1111111011110000",
    "1111111010111100",
    "1111111100101101",
    "1111111111000011",
    "1111111000110101",
    "1111110001001001",
    "1111101000100101",
    "1111011111110000",
    "1111010111001011",
    "1111001111010110",
    "1111001000100111",
    "1111000011010101",
    "1110111111110000",
    "1110111110000010",
    "1110111110001111",
    "1111000000010111",
    "1111000100011000",
    "1111001010010100",
    "1111010010001010",
    "1111011011111000",
    "1111100111011011",
    "1111110100101010",
    "1111111100110100",
    "1111101101110110",
    "1111011111101100",
    "1111010100000110",
    "1111001100110111",
    "1111001011101000",
    "1111010001001111",
    "1111011101010001",
    "1111101110000001",
    "1111111111010000",
    "1111101101101110",
    "1111100000000000",
    "1111010111101010",
    "1111010100111011",
    "1111010110111011",
    "1111011100000100",
    "1111100010111001",
    "1111101010010011",
    "1111110001110000",
    "1111111001000011",
    "1111111111111101",
    "1111111001110000",
    "1111110100111011",
    "1111110010000110",
    "1111110001101100",
    "1111110011100011",
    "1111110110111110",
    "1111111010110110",
    "1111111101111100",
    "1111111111001111",
    "1111111110000101",
    "1111111010010001",
    "1111110011111110",
    "1111101011100100",
    "1111100001100010",
    "1111010110100000",
    "1111001011000100",
    "1110111111110101",
    "1110110101010111",
    "1110101100000001",
    "1110100100000011",
    "1110011101100001",
    "1110011000011000",
    "1110010100100100",
    "1110010010000000",
    "1110010000101100",
    "1110010000101011",
    "1110010001110100",
    "1110010100001011",
    "1110010111101101",
    "1110011100101000",
    "1110100011001011",
    "1110101011101011",
    "1110110110010110",
    "1111000011001011",
    "1111010001110000",
    "1111100001001111",
    "1111110000100110",
    "1111111110101000",
    "1111110101101000",
    "1111101100111111",
    "1111100111101101",
    "1111100101101111",
    "1111100110110110",
    "1111101010110011",
    "1111110001011101",
    "1111111010110111",
    "1111111000100110",
    "1111101000110010",
    "1111010101111100",
    "1111000001001111",
    "1110101100101011",
    "1110011010101111",
    "1110001101100100",
    "1110000110011010",
    "1110000101000110",
    "1110001000011000",
    "1110001110011001",
    "1110010101011000",
    "1110011100001111",
    "1110100010101110",
    "1110101001000001",
    "1110101111100100",
    "1110110110011111",
    "1110111101101001",
    "1111000100101110",
    "1111001011010110",
    "1111010001100010",
    "1111010111100010",
    "1111011101110101",
    "1111100100111011",
    "1111101101000011",
    "1111110110000010",
    "1111111111011110",
    "1111110111000110",
    "1111101110001010",
    "1111100101111100",
    "1111011110101101",
    "1111011000100010",
    "1111010011100010",
    "1111001111111010",
    "1111001101110011",
    "1111001101100100",
    "1111001111100110",
    "1111010100010111",
    "1111011100001110",
    "1111100111010101",
    "1111110101011010",
    "1111111010010110",
    "1111101001010110",
    "1111011001001110",
    "1111001011100000",
    "1111000001011010",
    "1110111011100000",
    "1110111001101010",
    "1110111011001010",
    "1110111110111111",
    "1111000100000000",
    "1111001001011000",
    "1111001110011100",
    "1111010010111110",
    "1111010110111011",
    "1111011010011101",
    "1111011101111010",
    "1111100001100111",
    "1111100101111100",
    "1111101011000000",
    "1111110000111001",
    "1111110111011010",
    "1111111110000110",
    "1111111011101001",
    "1111110110101010",
    "1111110011100110",
    "1111110010110110",
    "1111110100011101",
    "1111110111111011",
    "1111111100010101",
    "1111111111011001",
    "1111111100011111",
    "1111111011110010",
    "1111111101111001",
    "1111111101000000",
    "1111110101010010",
    "1111101011110000",
    "1111100001110001",
    "1111011001000110",
    "1111010011011101",
    "1111010010001011",
    "1111010101110100",
    "1111011101111011",
    "1111101001010011",
    "1111110101111101",
    "1111111110001010",
    "1111110101001001",
    "1111110000100111",
    "1111110001100101",
    "1111111000001100",
    "1111111100001101",
    "1111101101010000",
    "1111011100111111",
    "1111001101100011",
    "1111000000110001",
    "1110110111101111",
    "1110110010101100",
    "1110110001001111",
    "1110110010100111",
    "1110110110000001",
    "1110111010111111",
    "1111000001011010",
    "1111001001010001",
    "1111010010100110",
    "1111011101001001",
    "1111101000100010",
    "1111110100010000",
    "1111111111110100",
    "1111110101000101",
    "1111101010101010",
    "1111100000111001",
    "1111010111110100",
    "1111001111011100",
    "1111000111111001",
    "1111000001001101",
    "1110111011100011",
    "1110110111000110",
    "1110110011111100",
    "1110110010001011",
    "1110110001110000",
    "1110110010011101",
    "1110110100000011",
    "1110110110001101",
    "1110111000101100",
    "1110111011011101",
    "1110111110101000",
    "1111000010011010",
    "1111000111000110",
    "1111001100111000",
    "1111010011110011",
    "1111011100000010",
    "1111100101111100",
    "1111110001101111",
    "1111111111010010",
    "1111110010001001",
    "1111100100000101",
    "1111010111111111",
    "1111001111001100",
    "1111001010000110",
    "1111001000000011",
    "1111000111100010",
    "1111000110101100",
    "1111000100000011",
    "1110111110111000",
    "1110110111100000",
    "1110101110111010",
    "1110100110100000",
    "1110011111101001",
    "1110011011001110",
    "1110011001101000",
    "1110011010101101",
    "1110011101111111",
    "1110100010111001",
    "1110101001000100",
    "1110110000001101",
    "1110111000010110",
    "1111000001011110",
    "1111001011100001",
    "1111010110010011",
    "1111100001010100",
    "1111101011101010",
    "1111110100011010",
    "1111111010101101",
    "1111111110000100",
    "1111111110011001",
    "1111111100000101",
    "1111110111101100",
    "1111110001111010",
    "1111101011010011",
    "1111100100010101",
    "1111011101010001",
    "1111010110010110",
    "1111001111110000",
    "1111001001101000",
    "1111000100010000",
    "1110111111111011",
    "1110111100111000",
    "1110111011011001",
    "1110111011011011",
    "1110111100110111",
    "1110111111011100",
    "1111000010111011",
    "1111000110111100",
    "1111001011010011",
    "1111001111110001",
    "1111010100010000",
    "1111011000101100",
    "1111011100111000",
    "1111100000100100",
    "1111100011001101",
    "1111100100001011",
    "1111100010110011",
    "1111011110101101",
    "1111010111110100",
    "1111001110101001",
    "1111000100010010",
    "1110111010000010",
    "1110110001011111",
    "1110101011111101",
    "1110101010011110",
    "1110101101100011",
    "1110110101000101",
    "1111000000000111",
    "1111001101001001",
    "1111011001111101",
    "1111100100010101",
    "1111101010001101",
    "1111101010001010",
    "1111100011101111",
    "1111010111101000",
    "1111000111101100",
    "1110110110011101",
    "1110100110111011",
    "1110011011100101",
    "1110010110001110",
    "1110010111011111",
    "1110011110111111",
    "1110101011101011",
    "1110111100010110",
    "1111001111110011",
    "1111100100111011",
    "1111111010100110",
    "1111110000100100",
    "1111011110000010",
    "1111001111000010",
    "1111000100001101",
    "1110111101011100",
    "1110111001111111",
    "1110111000100010",
    "1110110111110101",
    "1110110111000100",
    "1110110110000011",
    "1110110101001000",
    "1110110101000000",
    "1110110110010010",
    "1110111001010101",
    "1110111110001101",
    "1111000100110110",
    "1111001100111111",
    "1111010110011010",
    "1111100000111110",
    "1111101100011000",
    "1111111000001000",
    "1111111100100100",
    "1111110010101111",
    "1111101011001000",
    "1111100110001101",
    "1111100011111011",
    "1111100011110100",
    "1111100101001110",
    "1111100111011100",
    "1111101001111100",
    "1111101100100001",
    "1111101111001100",
    "1111110001111100",
    "1111110100101000",
    "1111110110111000",
    "1111111000001110",
    "1111111000001111",
    "1111110110101111",
    "1111110011111001",
    "1111110000001000",
    "1111101100000111",
    "1111101000100011",
    "1111100110000001",
    "1111100101000001",
    "1111100101111011",
    "1111101000111001",
    "1111101110000111",
    "1111110101011111",
    "1111111110110001",
    "1111110110100110",
    "1111101011101001",
    "1111100001101001",
    "1111011010000100",
    "1111010110010000",
    "1111010111001001",
    "1111011100111000",
    "1111100110110110",
    "1111110011110001",
    "1111111110000011",
    "1111110000011100",
    "1111100100111011",
    "1111011100100000",
    "1111010111101010",
    "1111010110011010",
    "1111011000011011",
    "1111011101010001",
    "1111100100100010",
    "1111101101111101",
    "1111111001010100",
    "1111111001101011",
    "1111101011101111",
    "1111011101101110",
    "1111010000110011",
    "1111000110000001",
    "1110111110001100",
    "1110111001101101",
    "1110111000011110",
    "1110111010000110",
    "1110111101111000",
    "1111000011001000",
    "1111001001001011",
    "1111001111011001",
    "1111010101001011",
    "1111011010000100",
    "1111011101101001",
    "1111011111101110",
    "1111100000010100",
    "1111011111101001",
    "1111011110001101",
    "1111011100100001",
    "1111011011000111",
    "1111011010011110",
    "1111011010111000",
    "1111011100100001",
    "1111011111010111",
    "1111100011001011",
    "1111100111101101",
    "1111101100101000",
    "1111110001110000",
    "1111110111000000",
    "1111111100011110",
    "1111111101110001",
    "1111110111111000",
    "1111110010001001",
    "1111101101000100",
    "1111101001001111",
    "1111100111001110",
    "1111100111010111",
    "1111101001110010",
    "1111101110011101",
    "1111110101011000",
    "1111111110100110",
    "1111110101101100",
    "1111100111011001",
    "1111010110111001",
    "1111000101011000",
    "1110110100111100",
    "1110101000010011",
    "1110100001111011",
    "1110100011100110",
    "1110101101110010",
    "1110111111011010",
    "1111010110000000",
    "1111101110000111",
    "1111111011101101",
    "1111101010010001",
    "1111011111001000",
    "1111011010011110",
    "1111011011011000",
    "1111100000001010",
    "1111100111000001",
    "1111101110011110",
    "1111110101011011",
    "1111111011010000",
    "1111111111100010",
    "1111111110000000",
    "1111111101100000",
    "1111111110110110",
    "1111111110010011",
    "1111111010101111",
    "1111110111011000",
    "1111110101001110",
    "1111110101010001",
    "1111111000001101",
    "1111111110010001",
    "1111111000101101",
    "1111101101011100",
    "1111100000110101",
    "1111010011111000",
    "1111000111100000",
    "1110111100011100",
    "1110110011000001",
    "1110101011001001",
    "1110100100011010",
    "1110011110010111",
    "1110011000101100",
    "1110010011010111",
    "1110001110101001",
    "1110001010111101",
    "1110001000110010",
    "1110001000011000",
    "1110001001110010",
    "1110001100111010",
    "1110010001100001",
    "1110010111011011",
    "1110011110101001",
    "1110100111011010",
    "1110110010000011",
    "1110111111000000",
    "1111001110011001",
    "1111011111111101",
    "1111110010101101",
    "1111111010110110",
    "1111101010100101",
    "1111011101111111",
    "1111010101110111",
    "1111010010001111",
    "1111010010010101",
    "1111010101000001",
    "1111011001010000",
    "1111011110011001",
    "1111100100011101",
    "1111101011110100",
    "1111110100101110",
    "1111111111000010",
    "1111110101111111",
    "1111101011101001",
    "1111100011011100",
    "1111011110101011",
    "1111011101111111",
    "1111100001010100",
    "1111100111110110",
    "1111110000010100",
    "1111111001010110",
    "1111111110010101",
    "1111110111110010",
    "1111110011100101",
    "1111110010000010",
    "1111110011001000",
    "1111110110100101",
    "1111111011110110",
    "1111111101101111",
    "1111110111000000",
    "1111110000101011",
    "1111101011010101",
    "1111100111011010",
    "1111100101001011",
    "1111100100110100",
    "1111100110011111",
    "1111101010010111",
    "1111110000011011",
    "1111111000011000",
    "1111111110011001",
    "1111110100111111",
    "1111101100100110",
    "1111100110010101",
    "1111100011000000",
    "1111100010110100",
    "1111100101101010",
    "1111101011000001",
    "1111110010001111",
    "1111111010101011",
    "1111111100001110",
    "1111110011001000",
    "1111101010100101",
    "1111100011001111",
    "1111011101100110",
    "1111011010001110",
    "1111011001010011",
    "1111011010111000",
    "1111011110110011",
    "1111100100101001",
    "1111101011111110",
    "1111110100010001",
    "1111111101000000",
    "1111111010010010",
    "1111110010001111",
    "1111101011010011",
    "1111100101110100",
    "1111100010000011",
    "1111100000000111",
    "1111100000000000",
    "1111100001110001",
    "1111100101011010",
    "1111101010111001",
    "1111110010000000",
    "1111111010010001",
    "1111111101000011",
    "1111110101000011",
    "1111101110110011",
    "1111101011010100",
    "1111101011011011",
    "1111101111101001",
    "1111111000010110",
    "1111111010011100",
    "1111101001100011",
    "1111010110100111",
    "1111000100000011",
    "1110110100100010",
    "1110101010011001",
    "1110100110111110",
    "1110101010010011",
    "1110110011010000",
    "1111000000000010",
    "1111001110101011",
    "1111011101010100",
    "1111101010011000",
    "1111110100010011",
    "1111111001101011",
    "1111111001011110",
    "1111110011001011",
    "1111100111001111",
    "1111010111001101",
    "1111000101011101",
    "1110110100101110",
    "1110100111011101",
    "1110011111011010",
    "1110011101010010",
    "1110100000111101",
    "1110101001110100",
    "1110110111000011",
    "1111000111101000",
    "1111011010010011",
    "1111101101011001",
    "1111111111001001",
    "1111110001111101",
    "1111100110111101",
    "1111011111110110",
    "1111011011111101",
    "1111011010000111",
    "1111011001001011",
    "1111011000011110",
    "1111010111111001",
    "1111010111100111",
    "1111011000001000",
    "1111011001101010",
    "1111011100001010",
    "1111011111010111",
    "1111100010110110",
    "1111100110011001",
    "1111101001111101",
    "1111101101110110",
    "1111110010011100",
    "1111111000001011",
    "1111111111011110",
    "1111110111001011",
    "1111101011010101",
    "1111011100110101",
    "1111001100001100",
    "1110111010101010",
    "1110101010000110",
    "1110011100011001",
    "1110010011000011",
    "1110001110101000",
    "1110001110110011",
    "1110010010100010",
    "1110011000100101",
    "1110011111110101",
    "1110100111100111",
    "1110101111011110",
    "1110110111000011",
    "1110111101111000",
    "1111000011011000",
    "1111000111000110",
    "1111001000110000",
    "1111001000101000",
    "1111000111011000",
    "1111000101111011",
    "1111000101001001",
    "1111000101100111",
    "1111000111011010",
    "1111001010011001",
    "1111001110010111",
    "1111010011001000",
    "1111011000110000",
    "1111011111010100",
    "1111100110110111",
    "1111101111001110",
    "1111111000000010",
    "1111111111001111",
    "1111110111010111",
    "1111110000110011",
    "1111101011111011",
    "1111101000110000",
    "1111100111000110",
    "1111100110100101",
    "1111100110110001",
    "1111100111001110",
    "1111100111100110",
    "1111100111101001",
    "1111100111001101",
    "1111100110001101",
    "1111100100101100",
    "1111100010101111",
    "1111100000011110",
    "1111011101111101",
    "1111011011010011",
    "1111011000101100",
    "1111010110011101",
    "1111010101000001",
    "1111010100111100",
    "1111010110101000",
    "1111011010010100",
    "1111011111111000",
    "1111100110110110",
    "1111101110100000",
    "1111110110001011",
    "1111111101010101",
    "1111111100001010",
    "1111110110001101",
    "1111110000100011",
    "1111101010111000",
    "1111100101001011",
    "1111011111100011",
    "1111011010011110",
    "1111010110011011",
    "1111010100000011",
    "1111010011101110",
    "1111010101101010",
    "1111011001111010",
    "1111100000001010",
    "1111100111110010",
    "1111101111110011",
    "1111110111000000",
    "1111111100001011",
    "1111111110001101",
    "1111111100011100",
    "1111110110101111",
    "1111101101110001",
    "1111100011000000",
    "1111011000011011",
    "1111010000010100",
    "1111001100100101",
    "1111001110101000",
    "1111010111000011",
    "1111100101011111",
    "1111111000110001",
    "1111110001000101",
    "1111011010101111",
    "1111000110110100",
    "1110110111101100",
    "1110101110111000",
    "1110101100110101",
    "1110110000111110",
    "1110111001111001",
    "1111000101110001",
    "1111010010111011",
    "1111011111111000",
    "1111101011100000",
    "1111110100111001",
    "1111111011010111",
    "1111111110101001",
    "1111111110110100",
    "1111111100011100",
    "1111111000011101",
    "1111110100001010",
    "1111110000110001",
    "1111101111010011",
    "1111110000001110",
    "1111110011011100",
    "1111111000011011",
    "1111111110011101",
    "1111111011001101",
    "1111110101010011",
    "1111110000001010",
    "1111101100000100",
    "1111101001001000",
    "1111100111011000",
    "1111100110111111",
    "1111101000001001",
    "1111101011000111",
    "1111110000000101",
    "1111110110111111",
    "1111111111011000",
    "1111110111110001",
    "1111101111111101",
    "1111101010110010",
    "1111101001101100",
    "1111101101101010",
    "1111110110110011",
    "1111111011101010",
    "1111101011100100",
    "1111011011000111",
    "1111001100101000",
    "1111000001111011",
    "1110111100000100",
    "1110111011001100",
    "1110111110110110",
    "1111000110001110",
    "1111010000100111",
    "1111011101100001",
    "1111101100011000",
    "1111111100011100",
    "1111110011100101",
    "1111100101011101",
    "1111011010110101",
    "1111010100111100",
    "1111010100000000",
    "1111010111010110",
    "1111011101100011",
    "1111100100111110",
    "1111101100001111",
    "1111110010100110",
    "1111110111110010",
    "1111111011110001",
    "1111111110100111",
    "1111111111110010",
    "1111111111101011",
    "1111111110101100",
    "1111111011011101",
    "1111110110110111",
    "1111110001100010",
    "1111101100010100",
    "1111100111111111",
    "1111100101010000",
    "1111100100011101",
    "1111100101110010",
    "1111101001001100",
    "1111101110011100",
    "1111110101001000",
    "1111111100110011",
    "1111111011001001",
    "1111110011011100",
    "1111101100101100",
    "1111100111100010",
    "1111100100011010",
    "1111100011100100",
    "1111100101000001",
    "1111101000100100",
    "1111101101101111",
    "1111110100000000",
    "1111111010101011",
    "1111111110110110",
    "1111111001001101",
    "1111110100101011",
    "1111110001011010",
    "1111101111010000",
    "1111101101111011",
    "1111101101000000",
    "1111101100000100",
    "1111101010110101",
    "1111101001000110",
    "1111100110110100",
    "1111100100000001",
    "1111100000111101",
    "1111011101110111",
    "1111011011000100",
    "1111011000110000",
    "1111010110111100",
    "1111010101010011",
    "1111010011010111",
    "1111010000101011",
    "1111001100111101",
    "1111001000011000",
    "1111000011011111",
    "1110111111010001",
    "1110111100101101",
    "1110111100110010",
    "1111000000001000",
    "1111000111000011",
    "1111010001100001",
    "1111011111010110",
    "1111101111111000",
    "1111111101111101",
    "1111101100000101",
    "1111011100110000",
    "1111010010010100",
    "1111001110011001",
    "1111010001100111",
    "1111011011001110",
    "1111101001010111",
    "1111111001110010",
    "1111110101101101",
    "1111100110110100",
    "1111011010011110",
    "1111010001001000",
    "1111001010110101",
    "1111000111100000",
    "1111000110110100",
    "1111001000001011",
    "1111001010101111",
    "1111001101010010",
    "1111001110110000",
    "1111001110001111",
    "1111001011100001",
    "1111000111000011",
    "1111000001110100",
    "1110111101000100",
    "1110111001111010",
    "1110111001010000",
    "1110111011100001",
    "1111000000111101",
    "1111001001011101",
    "1111010100100100",
    "1111100001011110",
    "1111101110111100",
    "1111111011101000",
    "1111111001110000",
    "1111110010001010",
    "1111101101111010",
    "1111101100110001",
    "1111101110001010",
    "1111110001100001",
    "1111110110100100",
    "1111111101011001",
    "1111111001101011",
    "1111101110101011",
    "1111100010000110",
    "1111010101001110",
    "1111001001111010",
    "1111000001111110",
    "1110111110101101",
    "1111000000100011",
    "1111000111000001",
    "1111010000111000",
    "1111011100100101",
    "1111101000100100",
    "1111110011010011",
    "1111111011011011",
    "1111111111110001",
    "1111111111100001",
    "1111111010011011",
    "1111110001001001",
    "1111100101001101",
    "1111011000110100",
    "1111001110011011",
    "1111001000001000",
    "1111000111001110",
    "1111001100000100",
    "1111010110001001",
    "1111100100100010",
    "1111110110000111",
    "1111110110001100",
    "1111100001110000",
    "1111001110000000",
    "1110111100100110",
    "1110101111000000",
    "1110100110001101",
    "1110100010100001",
    "1110100011011111",
    "1110101000001110",
    "1110101111110000",
    "1110111001011001",
    "1111000100110111",
    "1111010010000010",
    "1111100000100111",
    "1111101111111111",
    "1111111110111001",
    "1111110100001110",
    "1111101011000000",
    "1111100110011110",
    "1111100110110111",
    "1111101011011110",
    "1111110010111110",
    "1111111011101011",
    "1111111011111010",
    "1111110101000011",
    "1111110000011110",
    "1111101110011111",
    "1111101111000011",
    "1111110001110001",
    "1111110110000011",
    "1111111011001100",
    "1111111111100001",
    "1111111010110110",
    "1111110111010111",
    "1111110101010111",
    "1111110101000001",
    "1111110110010001",
    "1111111000111011",
    "1111111100101111",
    "1111111110100100",
    "1111111001011000",
    "1111110011111110",
    "1111101110101011",
    "1111101001101111",
    "1111100101011000",
    "1111100001110110",
    "1111011111010100",
    "1111011110000101",
    "1111011110100110",
    "1111100001011111",
    "1111100111011100",
    "1111110001000001",
    "1111111110001110",
    "1111110001100011",
    "1111011111111010",
    "1111001110101110",
    "1111000000000101",
    "1110110101100101",
    "1110110000000011",
    "1110101111011010",
    "1110110010111000",
    "1110111001000100",
    "1111000000100001",
    "1111000111111111",
    "1111001110011111",
    "1111010011101001",
    "1111010111101010",
    "1111011011011101",
    "1111100000000000",
    "1111100101111001",
    "1111101101000000",
    "1111110100011101",
    "1111111010111010",
    "1111111111001101",
    "1111111111001010",
    "1111111111110110",
    "1111111110011010",
    "1111111101010001",
    "1111111110000010",
    "1111111110101011",
    "1111111001001001",
    "1111110010001001",
    "1111101010111101",
    "1111100100110011",
    "1111100000101100",
    "1111011111011100",
    "1111100001010101",
    "1111100110011000",
    "1111101110001010",
    "1111110111111011",
    "1111111101010100",
    "1111110010110101",
    "1111101001101001",
    "1111100010100010",
    "1111011101110111",
    "1111011011011110",
    "1111011010111111",
    "1111011011110010",
    "1111011101010001",
    "1111011111000000",
    "1111100000101001",
    "1111100010000011",
    "1111100011010000",
    "1111100100011010",
    "1111100101110110",
    "1111101000000010",
    "1111101011100100",
    "1111110001000110",
    "1111111001001110",
    "1111111011101010",
    "1111101101100001",
    "1111011100011001",
    "1111001000111001",
    "1110110100000001",
    "1110011111100001",
    "1110001101001111",
    "1101111110111010",
    "1101110101100101",
    "1101110001100010",
    "1101110010000000",
    "1101110101101010",
    "1101111011000110",
    "1110000001011001",
    "1110001000010101",
    "1110010000001111",
    "1110011001100101",
    "1110100100011010",
    "1110101111111101",
    "1110111010101111",
    "1111000010110001",
    "1111000110010010",
    "1111000100001110",
    "1110111100110101",
    "1110110001011010",
    "1110100100000011",
    "1110010110111110",
    "1110001100001010",
    "1110000101000001",
    "1110000010010101",
    "1110000100011000",
    "1110001010111111",
    "1110010101110110",
    "1110100100001101",
    "1110110101000000",
    "1111000110100111",
    "1111010111000100",
    "1111100100011100",
    "1111101101001111",
    "1111110000110110",
    "1111101111101011",
    "1111101010111101",
    "1111100100010010",
    "1111011101001111",
    "1111010111001000",
    "1111010010101110",
    "1111010000100100",
    "1111010001001000",
    "1111010100101001",
    "1111011011010100",
    "1111100101000001",
    "1111110001010100",
    "1111111111011000",
    "1111110001110010",
    "1111100011011010",
    "1111010110011010",
    "1111001011100011",
    "1111000011010010",
    "1110111101111011",
    "1110111011101111",
    "1110111100111010",
    "1111000001101011",
    "1111001010000100",
    "1111010101110111",
    "1111100100100101",
    "1111110101011001",
    "1111111000111001",
    "1111100111101100",
    "1111011000001110",
    "1111001011011110",
    "1111000001110110",
    "1110111011011000",
    "1110110111100011",
    "1110110101101100",
    "1110110101000001",
    "1110110101000000",
    "1110110101010101",
    "1110110110000001",
    "1110110111010110",
    "1110111001110101",
    "1110111101111010",
    "1111000011111110",
    "1111001011111010",
    "1111010101001101",
    "1111011110111000",
    "1111100111101100",
    "1111101110011111",
    "1111110010100011",
    "1111110011110001",
    "1111110010111011",
    "1111110001010100",
    "1111110000100011",
    "1111110010000110",
    "1111110111000100",
    "1111111111111000",
    "1111110010100111",
    "1111100001101100",
    "1111001110011011",
    "1110111010111100",
    "1110101001111001",
    "1110011101110011",
    "1110011000100000",
    "1110011010101111",
    "1110100011111001",
    "1110110010011100",
    "1111000100100000",
    "1111011000011010",
    "1111101100110010",
    "1111111111011000",
    "1111101101001101",
    "1111011101110111",
    "1111010010011010",
    "1111001011101011",
    "1111001001110100",
    "1111001100000101",
    "1111010001001100",
    "1111010111011111",
    "1111011101101110",
    "1111100011010111",
    "1111101000100010",
    "1111101101111110",
    "1111110100011111",
    "1111111100100100",
    "1111111001101010",
    "1111101110101000",
    "1111100011000001",
    "1111010111101000",
    "1111001101010100",
    "1111000100100111",
    "1110111101111111",
    "1110111001011011",
    "1110110110110110",
    "1110110101110100",
    "1110110101110010",
    "1110110110011010",
    "1110110111011011",
    "1110111001000100",
    "1110111011110011",
    "1111000000010001",
    "1111000110111110",
    "1111010000000011",
    "1111011011000010",
    "1111100110111011",
    "1111110010010001",
    "1111111011101111",
    "1111111101100111",
    "1111111010001110",
    "1111111001111010",
    "1111111100000101",
    "1111111111111100",
    "1111111011011001",
    "1111110110110110",
    "1111110011010001",
    "1111110001010110",
    "1111110001101001",
    "1111110100001101",
    "1111111000101001",
    "1111111110000111",
    "1111111100100110",
    "1111111000101011",
    "1111110110111100",
    "1111110111110010",
    "1111111010111110",
    "1111111111111111",
    "1111111001111100",
    "1111110011100111",
    "1111101101100110",
    "1111101000010010",
    "1111100011111001",
    "1111100000100100",
    "1111011110010111",
    "1111011101010100",
    "1111011101010111",
    "1111011110100001",
    "1111100000101110",
    "1111100011111000",
    "1111100111110101",
    "1111101100100000",
    "1111110001101100",
    "1111110111001111",
    "1111111100110111",
    "1111111101101110",
    "1111111001000000",
    "1111110101010110",
    "1111110011000111",
    "1111110010011111",
    "1111110011011101",
    "1111110101110100",
    "1111111001001111",
    "1111111101011000",
    "1111111110000100",
    "1111111001010010",
    "1111110100001110",
    "1111101110101011",
    "1111101000010010",
    "1111100000100100",
    "1111010111001000",
    "1111001011110010",
    "1110111110110000",
    "1110110000110101",
    "1110100011000101",
    "1110010110101100",
    "1110001100100110",
    "1110000101010000",
    "1110000000100011",
    "1101111101111101",
    "1101111100110101",
    "1101111100101010",
    "1101111101000100",
    "1101111101111101",
    "1101111111010100",
    "1110000001001000",
    "1110000011010101",
    "1110000101110110",
    "1110001000100011",
    "1110001011100000",
    "1110001110110001",
    "1110010010100010",
    "1110010111000110",
    "1110011101001010",
    "1110100110000001",
    "1110110011000110",
    "1111000101010011",
    "1111011100001110",
    "1111110101110100",
    "1111110001010101",
    "1111011101001001",
    "1111010000100110",
    "1111001100111000",
    "1111010000111000",
    "1111011001111010",
    "1111100100111001",
    "1111101111010100",
    "1111110111111001",
    "1111111110100110",
    "1111111011111101",
    "1111110111001111",
    "1111110011000110",
    "1111101111111110",
    "1111101110011100",
    "1111101110111000",
    "1111110001000010",
    "1111110100000101",
    "1111110110111010",
    "1111111000100100",
    "1111111000100011",
    "1111110110111011",
    "1111110100000100",
    "1111110000011111",
    "1111101100101011",
    "1111101000111011",
    "1111100101011111",
    "1111100010011001",
    "1111011111110000",
    "1111011101100100",
    "1111011011110111",
    "1111011010011110",
    "1111011001011011",
    "1111011000101100",
    "1111011000010000",
    "1111011000001110",
    "1111011000101100",
    "1111011001101000",
    "1111011010111101",
    "1111011100011011",
    "1111011101110010",
    "1111011110110000",
    "1111011111011001",
    "1111011111110110",
    "1111100000100100",
    "1111100010000000",
    "1111100100100100",
    "1111101000101101",
    "1111101110101011",
    "1111110110110000",
    "1111111110111101",
    "1111110010101100",
    "1111100101000110",
    "1111010111011010",
    "1111001011001010",
    "1111000001111101",
    "1110111100110101",
    "1110111100001100",
    "1110111111011110",
    "1111000101010111",
    "1111001100001100",
    "1111010010010000",
    "1111010110010010",
    "1111010111100010",
    "1111010101110110",
    "1111010001100110",
    "1111001011011001",
    "1111000100000000",
    "1110111100000111",
    "1110110100011010",
    "1110101101011100",
    "1110100111101101",
    "1110100011100100",
    "1110100001001100",
    "1110100000100110",
    "1110100001101001",
    "1110100100000101",
    "1110100111101111",
    "1110101100100000",
    "1110110010010111",
    "1110111001011110",
    "1111000001111000",
    "1111001011100000",
    "1111010110001001",
    "1111100001010111",
    "1111101100100110",
    "1111110111001000",
    "1111111111100100",
    "1111110111111111",
    "1111110010010001",
    "1111101110011110",
    "1111101100011111",
    "1111101100001000",
    "1111101101001010",
    "1111101111010011",
    "1111110010001100",
    "1111110101011011",
    "1111111000101010",
    "1111111011100011",
    "1111111101111001",
    "1111111111100111",
    "1111111111001000",
    "1111111110001111",
    "1111111101010111",
    "1111111100001101",
    "1111111010100101",
    "1111111000011011",
    "1111110101110010",
    "1111110010110010",
    "1111101111100011",
    "1111101100001101",
    "1111101000101100",
    "1111100100110100",
    "1111100000010010",
    "1111011010110111",
    "1111010100100100",
    "1111001101110011",
    "1111000111100111",
    "1111000011010010",
    "1111000010010100",
    "1111000101110100",
    "1111001110001001",
    "1111011010011110",
    "1111101001000110",
    "1111110111100110",
    "1111111100011010",
    "1111110100110110",
    "1111110010101001",
    "1111110101110001",
    "1111111101101101",
    "1111110110001010",
    "1111100110010101",
    "1111010011010011",
    "1110111110010001",
    "1110101001001011",
    "1110010110100101",
    "1110001001000100",
    "1110000010010000",
    "1110000010100001",
    "1110001000100011",
    "1110010010001011",
    "1110011100111111",
    "1110100111001011",
    "1110101111111111",
    "1110110111011011",
    "1110111110000000",
    "1111000100001010",
    "1111001001111100",
    "1111001111001101",
    "1111010011101110",
    "1111010111011111",
    "1111011010111010",
    "1111011110101011",
    "1111100011011000",
    "1111101001010101",
    "1111110000010101",
    "1111110111110011",
    "1111111111000111",
    "1111111010001010",
    "1111110100011001",
    "1111101111100111",
    "1111101011101111",
    "1111101000100111",
    "1111100110000110",
    "1111100011111110",
    "1111100010000110",
    "1111100000010100",
    "1111011110100100",
    "1111011100110101",
    "1111011011010100",
    "1111011010001110",
    "1111011001110101",
    "1111011010001111",
    "1111011011011001",
    "1111011101000101",
    "1111011111000111",
    "1111100001010000",
    "1111100011110001",
    "1111100110111100",
    "1111101011011001",
    "1111110001101100",
    "1111111010011011",
    "1111111010000111",
    "1111101100010000",
    "1111011100111010",
    "1111001101110000",
    "1111000000110001",
    "1110110111110101",
    "1110110100001011",
    "1110110110001011",
    "1110111101010010",
    "1111001000011101",
    "1111010110011010",
    "1111100110000100",
    "1111110110010111",
    "1111111001110010",
    "1111101011110000",
    "1111100000111000",
    "1111011010001111",
    "1111011000011010",
    "1111011011000010",
    "1111100001001000",
    "1111101001001011",
    "1111110001101011",
    "1111111001011110",
    "1111111111111000",
    "1111111011010100",
    "1111111000011000",
    "1111110111011001",
    "1111111000101011",
    "1111111100011000",
    "1111111101100011",
    "1111110101100111",
    "1111101100100100",
    "1111100011010000",
    "1111011010011110",
    "1111010010101110",
    "1111001100010100",
    "1111000111011010",
    "1111000100001011",
    "1111000011000000",
    "1111000100001010",
    "1111000111110001",
    "1111001101101000",
    "1111010101000101",
    "1111011101000111",
    "1111100100100000",
    "1111101010001100",
    "1111101101010100",
    "1111101101100110",
    "1111101011001000",
    "1111100110010101",
    "1111011111111010",
    "1111011000100111",
    "1111010001010000",
    "1111001010110000",
    "1111000101111011",
    "1111000011011100",
    "1111000011111001",
    "1111000111100101",
    "1111001110101001",
    "1111011001000100",
    "1111100110100111",
    "1111110110110101",
    "1111110111000001",
    "1111100100001101",
    "1111010010001010",
    "1111000010010010",
    "1110110101110001",
    "1110101101000101",
    "1110101000010000",
    "1110100110101111",
    "1110100111111110",
    "1110101011101000",
    "1110110001110100",
    "1110111011000111",
    "1111001000001100",
    "1111011001000111",
    "1111101100111010",
    "1111111110101101",
    "1111101100111101",
    "1111100000111011",
    "1111011100101101",
    "1111100000111000",
    "1111101100010110",
    "1111111100111001",
    "1111110000001011",
    "1111011101100110",
    "1111001101101000",
    "1111000010001000",
    "1110111100011100",
    "1110111101011001",
    "1111000101000001",
    "1111010010100100",
    "1111100100010000",
    "1111110111100010",
    "1111110110011011",
    "1111101000011001",
    "1111100000001100",
    "1111011110101000",
    "1111100011011101",
    "1111101101100000",
    "1111111010111110",
    "1111110110001010",
    "1111100111111010",
    "1111011011111101",
    "1111010011011100",
    "1111001110110110",
    "1111001110000000",
    "1111010000001000",
    "1111010100001010",
    "1111011001000110",
    "1111011110010111",
    "1111100011101111",
    "1111101001010011",
    "1111101111001011",
    "1111110101011110",
    "1111111100000110",
    "1111111101001011",
    "1111110110111011",
    "1111110001100000",
    "1111101101010110",
    "1111101010100111",
    "1111101001010101",
    "1111101001011001",
    "1111101010100000",
    "1111101100010001",
    "1111101110001011",
    "1111101111100111",
    "1111110000000110",
    "1111101111010111",
    "1111101101011111",
    "1111101011000010",
    "1111101000110110",
    "1111100111110110",
    "1111101000110101",
    "1111101100000100",
    "1111110001010101",
    "1111110111110111",
    "1111111110011110",
    "1111111100000101",
    "1111111001000111",
    "1111111001011100",
    "1111111101100100",
    "1111111010011101",
    "1111101111010101",
    "1111100010001010",
    "1111010100100111",
    "1111001000011110",
    "1110111111010110",
    "1110111010010110",
    "1110111010000001",
    "1110111110010001",
    "1111000110101101",
    "1111010010100110",
    "1111100000110110",
    "1111110000000110",
    "1111111110101001",
    "1111110101000010",
    "1111101100001100",
    "1111100111001101",
    "1111100101101110",
    "1111100110101011",
    "1111101000110111",
    "1111101011010010",
    "1111101101011101",
    "1111101111011100",
    "1111110001100011",
    "1111110100000010",
    "1111110110110011",
    "1111111001011000",
    "1111111011001001",
    "1111111011100001",
    "1111111010010011",
    "1111110111101111",
    "1111110100011110",
    "1111110001010010",
    "1111101110111011",
    "1111101110000001",
    "1111101111000010",
    "1111110010011001",
    "1111111000100100",
    "1111111101111111",
    "1111110001000000",
    "1111100000011111",
    "1111001101000101",
    "1110111000001001",
    "1110100011100010",
    "1110010001001111",
    "1110000010111001",
    "1101111001100111",
    "1101110101100100",
    "1101110110010110",
    "1101111011010001",
    "1110000011100010",
    "1110001110011110",
    "1110011011101111",
    "1110101010111101",
    "1110111011110111",
    "1111001101110101",
    "1111011111111101",
    "1111110001000010",
    "1111111111111000",
    "1111110100011101",
    "1111101100011110",
    "1111101000000001",
    "1111100110100100",
    "1111100111010000",
    "1111101001010101",
    "1111101100010100",
    "1111101111111011",
    "1111110100000110",
    "1111111000101011",
    "1111111101001010",
    "1111111111001011",
    "1111111101011111",
    "1111111110101010",
    "1111111100110100",
    "1111110101011001",
    "1111101100001110",
    "1111100011001011",
    "1111011100010001",
    "1111011001010000",
    "1111011011010001",
    "1111100010101011",
    "1111101111000101",
    "1111111111100100",
    "1111101101011010",
    "1111011001110111",
    "1111000111111111",
    "1110111001111111",
    "1110110001100110",
    "1110101111110101",
    "1110110100101001",
    "1110111111001100",
    "1111001101110010",
    "1111011110010010",
    "1111101110100100",
    "1111111100101000",
    "1111111000111111",
    "1111110011001111",
    "1111110010011010",
    "1111110110001110",
    "1111111101111101",
    "1111110111011110",
    "1111101011011001",
    "1111011111000100",
    "1111010011100001",
    "1111001001100011",
    "1111000001100001",
    "1110111011011001",
    "1110110110111001",
    "1110110011101001",
    "1110110001001111",
    "1110101111010100",
    "1110101101110000",
    "1110101100011011",
    "1110101011011001",
    "1110101010110101",
    "1110101011000001",
    "1110101100000101",
    "1110101110010001",
    "1110110001011010",
    "1110110101011111",
    "1110111010001111",
    "1110111111101001",
    "1111000101110111",
    "1111001101010100",
    "1111010110101100",
    "1111100010100111",
    "1111110001010101",
    "1111111101100111",
    "1111101011100000",
    "1111011010000100",
    "1111001011000010",
    "1110111111110110",
    "1110111001001100",
    "1110110110111111",
    "1110111000101101",
    "1110111101100001",
    "1111000100101010",
    "1111001101010110",
    "1111010110101100",
    "1111011111100110",
    "1111100110111000",
    "1111101011010101",
    "1111101100001110",
    "1111101001011111",
    "1111100011111001",
    "1111011101000100",
    "1111010111000011",
    "1111010011110110",
    "1111010101000001",
    "1111011011010001",
    "1111100110011100",
    "1111110101011001",
    "1111111001101001",
    "1111101000111010",
    "1111011010011000",
    "1111001111010100",
    "1111001000010000",
    "1111000100101111",
    "1111000011111000",
    "1111000100100101",
    "1111000110001000",
    "1111001000000100",
    "1111001010100011",
    "1111001101110000",
    "1111010001111110",
    "1111010111010000",
    "1111011101011100",
    "1111100100001101",
    "1111101011000001",
    "1111110001011100",
    "1111110110111101",
    "1111111011001101",
    "1111111101110110",
    "1111111110110010",
    "1111111110000101",
    "1111111100000110",
    "1111111001100001",
    "1111110111001101",
    "1111110101111111",
    "1111110110011110",
    "1111111000111011",
    "1111111101010001",
    "1111111100110100",
    "1111110101111101",
    "1111101110110001",
    "1111100111111110",
    "1111100010001101",
    "1111011110000101",
    "1111011011111010",
    "1111011011101010",
    "1111011101000000",
    "1111011111010001",
    "1111100001100111",
    "1111100011010011",
    "1111100011110100",
    "1111100010111110",
    "1111100000110110",
    "1111011101110010",
    "1111011010000100",
    "1111010110000001",
    "1111010001101001",
    "1111001100110101",
    "1111000111010000",
    "1111000000010111",
    "1110110111100011",
    "1110101100010011",
    "1110011110011110",
    "1110001110110000",
    "1101111110011110",
    "1101101111100011",
    "1101100100000000",
    "1101011101100001",
    "1101011101000000",
    "1101100010100001",
    "1101101101010111",
    "1101111100100110",
    "1110001111000000",
    "1110100011011101",
    "1110111000100000",
    "1111001100100001",
    "1111011101101101",
    "1111101010011001",
    "1111110001010111",
    "1111110010010110",
    "1111101110000100",
    "1111100110010010",
    "1111011101000101",
    "1111010100101010",
    "1111001110100011",
    "1111001011011110",
    "1111001011011011",
    "1111001101101110",
    "1111010001010010",
    "1111010100111011",
    "1111010111101000",
    "1111011000101111",
    "1111010111110111",
    "1111010101001000",
    "1111010000111011",
    "1111001011111000",
    "1111000110101111",
    "1111000010001000",
    "1110111110100110",
    "1110111100011110",
    "1110111100000001",
    "1110111101010010",
    "1111000000010100",
    "1111000101000000",
    "1111001011000010",
    "1111010010000101",
    "1111011001101011",
    "1111100001011001",
    "1111101000110010",
    "1111101111101010",
    "1111110101110100",
    "1111111011000100",
    "1111111111001100",
    "1111111110001101",
    "1111111101110100",
    "1111111111101101",
    "1111111010000110",
    "1111110001100000",
    "1111100110111011",
    "1111011011111010",
    "1111010010011001",
    "1111001011111000",
    "1111001001011001",
    "1111001010111101",
    "1111001111111101",
    "1111010111010101",
    "1111011111111000",
    "1111101000011111",
    "1111110000000101",
    "1111110101100101",
    "1111110111111111",
    "1111110110011010",
    "1111110000011000",
    "1111100110000011",
    "1111011000100000",
    "1111001001011101",
    "1110111011000010",
    "1110101111001010",
    "1110100111001011",
    "1110100011100100",
    "1110100011111011",
    "1110100111011011",
    "1110101101001010",
    "1110110100011100",
    "1110111100111101",
    "1111000110110001",
    "1111010010000000",
    "1111011110101011",
    "1111101100100001",
    "1111111011000001",
    "1111110110100100",
    "1111101001000101",
    "1111011101001100",
    "1111010011010111",
    "1111001011110000",
    "1111000110010110",
    "1111000010111110",
    "1111000001010111",
    "1111000001010010",
    "1111000010011111",
    "1111000100110100",
    "1111001000001011",
    "1111001100011110",
    "1111010001101100",
    "1111010111110101",
    "1111011110111010",
    "1111100110110000",
    "1111101111000101",
    "1111110111011111",
    "1111111111011011",
    "1111111001100010",
    "1111110011110110",
    "1111101111100101",
    "1111101100101101",
    "1111101011000011",
    "1111101010011101",
    "1111101010110101",
    "1111101100001010",
    "1111101110011010",
    "1111110001100101",
    "1111110101100010",
    "1111111010000111",
    "1111111111010000",
    "1111111011000010",
    "1111110100100110",
    "1111101100111001",
    "1111100011010000",
    "1111010111001001",
    "1111001000100010",
    "1110111000001011",
    "1110100111100101",
    "1110011000100111",
    "1110001100111000",
    "1110000101011111",
    "1110000010100001",
    "1110000011011010",
    "1110000111001110",
    "1110001101001100",
    "1110010101001000",
    "1110011111011001",
    "1110101100011100",
    "1110111100010001",
    "1111001101111101",
    "1111011111110000",
    "1111101111011110",
    "1111111011001011",
    "1111111110001100",
    "1111111100100111",
    "1111111110101110",
    "1111111101010000",
    "1111111001001100",
    "1111110110010001",
    "1111110100111101",
    "1111110101000110",
    "1111110110001000",
    "1111110111011000",
    "1111111000010010",
    "1111111000100001",
    "1111110111111101",
    "1111110110100101",
    "1111110100100000",
    "1111110001111001",
    "1111101110111110",
    "1111101100000111",
    "1111101001101010",
    "1111100111110111",
    "1111100110110010",
    "1111100110010011",
    "1111100110001000",
    "1111100101110110",
    "1111100101000101",
    "1111100011100010",
    "1111100000111101",
    "1111011101001111",
    "1111011000011000",
    "1111010010011100",
    "1111001011100101",
    "1111000100010101",
    "1110111101011100",
    "1110110111111001",
    "1110110100110011",
    "1110110100111011",
    "1110111000101101",
    "1110111111111000",
    "1111001001101101",
    "1111010101001011",
    "1111100001011001",
    "1111101101101010",
    "1111111001011111",
    "1111111011100100",
    "1111110010001100",
    "1111101011001011",
    "1111100111011011",
    "1111100111101001",
    "1111101100000111",
    "1111110100110000",
    "1111111110110110",
    "1111101111011000",
    "1111011101100001",
    "1111001010010011",
    "1110110111000100",
    "1110100101100100",
    "1110010111100000",
    "1110001110010111",
    "1110001010110111",
    "1110001100110011",
    "1110010011001000",
    "1110011100011001",
    "1110100111000110",
    "1110110010001000",
    "1110111100110111",
    "1111000110111111",
    "1111010000011010",
    "1111011000111110",
    "1111100000010010",
    "1111100101111001",
    "1111101001011011",
    "1111101010101111",
    "1111101010001101",
    "1111101000100100",
    "1111100110111100",
    "1111100110011110",
    "1111101000001010",
    "1111101100100011",
    "1111110011100110",
    "1111111100100100",
    "1111111001101001",
    "1111110000100001",
    "1111101001001100",
    "1111100100011111",
    "1111100010101011",
    "1111100011100111",
    "1111100111000010",
    "1111101100101101",
    "1111110100101100",
    "1111111111010010",
    "1111110011001101",
    "1111100010111011",
    "1111010000100100",
    "1110111101101101",
    "1110101100010100",
    "1110011110010110",
    "1110010101001000",
    "1110010001000011",
    "1110010001100001",
    "1110010101010010",
    "1110011011000010",
    "1110100001110001",
    "1110101001000111",
    "1110110001000111",
    "1110111010000111",
    "1111000100011111",
    "1111010000011111",
    "1111011110001100",
    "1111101101011000",
    "1111111101101100",
    "1111110001100010",
    "1111100001011110",
    "1111010011011000",
    "1111001000110000",
    "1111000010101100",
    "1111000001110110",
    "1111000110001110",
    "1111001111000101",
    "1111011011000001",
    "1111101000000110",
    "1111110100001101",
    "1111111101011110",
    "1111111101100010",
    "1111111101101000",
    "1111111101001000",
    "1111110011010100",
    "1111100101110100",
    "1111010101111110",
    "1111000101100101",
    "1110110110101010",
    "1110101011001001",
    "1110100100100010",
    "1110100011100100",
    "1110100111111110",
    "1110110000101011",
    "1110111100000111",
    "1111001000110000",
    "1111010101010101",
    "1111100000111001",
    "1111101010110011",
    "1111110010011101",
    "1111110111011100",
    "1111111001011110",
    "1111111000011101",
    "1111110100101011",
    "1111101110101111",
    "1111100111011000",
    "1111011111011001",
    "1111010111010011",
    "1111001111011110",
    "1111001000001001",
    "1111000001101100",
    "1110111100101011",
    "1110111001110100",
    "1110111001110000",
    "1110111100110111",
    "1111000011000110",
    "1111001100001001",
    "1111010111010101",
    "1111100100000110",
    "1111110001110011",
    "1111111111110111",
    "1111110010010101",
    "1111100101101100",
    "1111011011000010",
    "1111010011010000",
    "1111001110111000",
    "1111001110000100",
    "1111010000011001",
    "1111010101001000",
    "1111011011010100",
    "1111100010001111",
    "1111101001011011",
    "1111110000111011",
    "1111111000111111",
    "1111111110000110",
    "1111110100010000",
    "1111101001100000",
    "1111011110001100",
    "1111010010111001",
    "1111001000011010",
    "1110111111100110",
    "1110111001010001",
    "1110110110000001",
    "1110110110000001",
    "1110111000111111",
    "1110111110010001",
    "1111000100110110",
    "1111001011110010",
    "1111010010000101",
    "1111010111001110",
    "1111011010111000",
    "1111011101000100",
    "1111011101111111",
    "1111011110000100",
    "1111011101110011",
    "1111011101111011",
    "1111011111001000",
    "1111100010001000",
    "1111100111010111",
    "1111101110111101",
    "1111111000100101",
    "1111111100100010",
    "1111110001100111",
    "1111100111101101",
    "1111011111110101",
    "1111011010100011",
    "1111010111111110",
    "1111010111101100",
    "1111011001001001",
    "1111011011101111",
    "1111011111000101",
    "1111100011001011",
    "1111101000011010",
    "1111101111011001",
    "1111111000110000",
    "1111111011001001",
    "1111101100101100",
    "1111011100111100",
    "1111001101100001",
    "1111000000011001",
    "1110110111001000",
    "1110110010110001",
    "1110110011100110",
    "1110111000111110",
    "1111000001111000",
    "1111001101000100",
    "1111011001011000",
    "1111100101111100",
    "1111110010000111",
    "1111111101011000",
    "1111111000101000",
    "1111110000011011",
    "1111101010010100",
    "1111100110101000",
    "1111100101011111",
    "1111100110101101",
    "1111101010000000",
    "1111101111000101",
    "1111110101101110",
    "1111111101111010",
    "1111111000010100",
    "1111101101010111",
    "1111100001110110",
    "1111010110110110",
    "1111001101100110",
    "1111000111010001",
    "1111000100101110",
    "1111000110010110",
    "1111001100010001",
    "1111010110001000",
    "1111100011001111",
    "1111110010001111",
    "1111111110101111",
    "1111110010001011",
    "1111101010010001",
    "1111101000101011",
    "1111101101111110",
    "1111111001101000",
    "1111110101110100",
    "1111100010011100",
    "1111001110100001",
    "1110111100010100",
    "1110101101111111",
    "1110100101010011",
    "1110100011101001",
    "1110101001100111",
    "1110110111000011",
    "1111001010101111",
    "1111100010010101",
    "1111111010111110",
    "1111101110011011",
    "1111011100011011",
    "1111010000011010",
    "1111001010101101",
    "1111001010011110",
    "1111001110010100",
    "1111010100111001",
    "1111011101001001",
    "1111100110010110",
    "1111110000001011",
    "1111111010001111",
    "1111111011111001",
    "1111110010111111",
    "1111101011101111",
    "1111100110111000",
    "1111100100111001",
    "1111100101111001",
    "1111101001101011",
    "1111101111101100",
    "1111110111001110",
    "1111111111100110",
    "1111110111111000",
    "1111101111111101",
    "1111101001010000",
    "1111100100011000",
    "1111100001110000",
    "1111100001011111",
    "1111100011100110",
    "1111100111101100",
    "1111101101010001",
    "1111110011101001",
    "1111111010000000",
    "1111111111100000",
    "1111111100100110",
    "1111111010111010",
    "1111111011100111",
    "1111111110011111",
    "1111111100111111",
    "1111110111110011",
    "1111110010110101",
    "1111101110111101",
    "1111101100110010",
    "1111101100011010",
    "1111101101100011",
    "1111101111011100",
    "1111110001010001",
    "1111110010001110",
    "1111110001110110",
    "1111110000000111",
    "1111101101011101",
    "1111101010101110",
    "1111101000110110",
    "1111101000101100",
    "1111101010101110",
    "1111101111000101",
    "1111110101011100",
    "1111111101010011",
    "1111111001110000",
    "1111110000001110",
    "1111100110010010",
    "1111011100010001",
    "1111010010100110",
    "1111001001111001",
    "1111000010110110",
    "1110111101111101",
    "1110111011011011",
    "1110111011000010",
    "1110111100010100",
    "1110111110110000",
    "1111000010000011",
    "1111000110001011",
    "1111001011010001",
    "1111010001100001",
    "1111011000101101",
    "1111100000010100",
    "1111100111010110",
    "1111101100110011",
    "1111101111110100",
    "1111110000000001",
    "1111101101101000",
    "1111101001011000",
    "1111100100001011",
    "1111011111000000",
    "1111011010100011",
    "1111010111010110",
    "1111010101101001",
    "1111010101011011",
    "1111010110101100",
    "1111011001001110",
    "1111011100101110",
    "1111100000111001",
    "1111100101011000",
    "1111101001110110",
    "1111101110000011",
    "1111110001110010",
    "1111110100111001",
    "1111110111010000",
    "1111111000110110",
    "1111111001101011",
    "1111111001111000",
    "1111111001100111",
    "1111111001000011",
    "1111111000010011",
    "1111110111011000",
    "1111110110001110",
    "1111110100110010",
    "1111110011000010",
    "1111110001001101",
    "1111101111101011",
    "1111101110111100",
    "1111101111100011",
    "1111110001111101",
    "1111110110011111",
    "1111111101010000",
    "1111111001110101",
    "1111101111010110",
    "1111100100001011",
    "1111011001101111",
    "1111010001110011",
    "1111001110001001",
    "1111010000001010",
    "1111011000010001",
    "1111100101110001",
    "1111110110100100",
    "1111111000000111",
    "1111101001010100",
    "1111011111011001",
    "1111011011101011",
    "1111011110010001",
    "1111100110001101",
    "1111110001111010",
    "1111111111101011",
    "1111110010000011",
    "1111100100101100",
    "1111011001011000",
    "1111010001000101",
    "1111001100100000",
    "1111001100000010",
    "1111001111011100",
    "1111010101111100",
    "1111011110001111",
    "1111100110110001",
    "1111101110000111",
    "1111110011010000",
    "1111110101110001",
    "1111110101110111",
    "1111110100000001",
    "1111110000111010",
    "1111101101001000",
    "1111101001000010",
    "1111100100110011",
    "1111100000010111",
    "1111011011101101",
    "1111010110101101",
    "1111010001011010",
    "1111001011110101",
    "1111000110000110",
    "1111000000011010",
    "1110111010111100",
    "1110110101111001",
    "1110110001011100",
    "1110101101101001",
    "1110101010100000",
    "1110100111110111",
    "1110100101011111",
    "1110100011000110",
    "1110100000011010",
    "1110011101001110",
    "1110011001100010",
    "1110010101100100",
    "1110010001110100",
    "1110001110111111",
    "1110001101110101",
    "1110001111001100",
    "1110010011100100",
    "1110011011001001",
    "1110100101100100",
    "1110110001110100",
    "1110111110011110",
    "1111001001110101",
    "1111010010010111",
    "1111010110111001",
    "1111010111000110",
    "1111010011011000",
    "1111001100111100",
    "1111000101011111",
    "1110111111000000",
    "1110111011011001",
    "1110111100000111",
    "1111000010000110",
    "1111001101101000",
    "1111011110000000",
    "1111110001110010",
    "1111111001001010",
    "1111100101010101",
    "1111010100110011",
    "1111001000111010",
    "1111000010000000",
    "1110111111011010",
    "1110111111110110",
    "1111000001110000",
    "1111000011111110",
    "1111000101110100",
    "1111000111011011",
    "1111001001101010",
    "1111001101111101",
    "1111010101110100",
    "1111100010010100",
    "1111110011010000",
    "1111111000101110",
    "1111100100000110",
    "1111010001110000",
    "1111000100000001",
    "1110111100010110",
    "1110111010101101",
    "1110111101111010",
    "1111000011111110",
    "1111001010110111",
    "1111010000110000",
    "1111010100011101",
    "1111010101100000",
    "1111010011111011",
    "1111010000000101",
    "1111001010100011",
    "1111000100000101",
    "1110111101100000",
    "1110110111101100",
    "1110110011100100",
    "1110110001110110",
    "1110110010111000",
    "1110110110101000",
    "1110111100101011",
    "1111000100011000",
    "1111001101000010",
    "1111010110000011",
    "1111011111001101",
    "1111101000101100",
    "1111110010111010",
    "1111111110010111",
    "1111110100110110",
    "1111100111011010",
    "1111011010011011",
    "1111001111011010",
    "1111000111110001",
    "1111000100100000",
    "1111000110000001",
    "1111001100001001",
    "1111010110010010",
    "1111100011011100",
    "1111110010001100",
    "1111111111001101",
    "1111110011000001",
    "1111101011011101",
    "1111101010100000",
    "1111110001010101",
    "1111111111110110",
    "1111101011100110",
    "1111010100000011",
    "1110111101001010",
    "1110101010010100",
    "1110011101111011",
    "1110011000111001",
    "1110011010100011",
    "1110100001011001",
    "1110101011100101",
    "1110110111101010",
    "1111000100101111",
    "1111010010010111",
    "1111100000010100",
    "1111101110001010",
    "1111111011001011",
    "1111111001011100",
    "1111110000100100",
    "1111101010100101",
    "1111100111011001",
    "1111100110010101",
    "1111100110011101",
    "1111100110110011",
    "1111100110101101",
    "1111100101110001",
    "1111100011111000",
    "1111100001001100",
    "1111011101110111",
    "1111011010000001",
    "1111010101110110",
    "1111010001010101",
    "1111001100100101",
    "1111000111101010",
    "1111000010110001",
    "1110111110001100",
    "1110111010010100",
    "1110110111101100",
    "1110110110101100",
    "1110110111101101",
    "1110111010111010",
    "1111000000000111",
    "1111000110111100",
    "1111001110110000",
    "1111010110110110",
    "1111011110100100",
    "1111100101011011",
    "1111101011001111",
    "1111110000000000",
    "1111110100000101",
    "1111111000001010",
    "1111111101010110",
    "1111111011000100",
    "1111110000001000",
    "1111100001011100",
    "1111001111101000",
    "1110111100010110",
    "1110101010010001",
    "1110011100001100",
    "1110010100011000",
    "1110010011111011",
    "1110011010101010",
    "1110100111011101",
    "1110111000100011",
    "1111001011110101",
    "1111011111001010",
    "1111110000011111",
    "1111111110001000",
    "1111111001000010",
    "1111110101100000",
    "1111110110110101",
    "1111111100000000",
    "1111111100010001",
    "1111110011000111",
    "1111101000111100",
    "1111011101101001",
    "1111010000111110",
    "1111000011000001",
    "1110110100101001",
    "1110100111001101",
    "1110011100011011",
    "1110010101101100",
    "1110010011101111",
    "1110010110010110",
    "1110011100100101",
    "1110100101000000",
    "1110101110001001",
    "1110110110101010",
    "1110111101011100",
    "1111000001100100",
    "1111000010100001",
    "1111000000001010",
    "1110111010110111",
    "1110110011100110",
    "1110101011100011",
    "1110100100001011",
    "1110011110110000",
    "1110011100001001",
    "1110011100110111",
    "1110100000111101",
    "1110101000010001",
    "1110110010011100",
    "1110111110111101",
    "1111001101000000",
    "1111011011100011",
    "1111101001010011",
    "1111110100111011",
    "1111111101010000",
    "1111111110011010",
    "1111111110011000",
    "1111111101101011",
    "1111110110100011",
    "1111101101000011",
    "1111100001111101",
    "1111010101110111",
    "1111001001010110",
    "1110111100110011",
    "1110110000110001",
    "1110100101110010",
    "1110011100100110",
    "1110010101110100",
    "1110010010000010",
    "1110010001101110",
    "1110010101001110",
    "1110011101000010",
    "1110101001100111",
    "1110111011000111",
    "1111010001000101",
    "1111101001101100",
    "1111111101110001",
    "1111101000100110",
    "1111011001011110",
    "1111010001110100",
    "1111010001011010",
    "1111010110011101",
    "1111011110101000",
    "1111100111101100",
    "1111110000011000",
    "1111111000010001",
    "1111111111100001",
    "1111111001110010",
    "1111110100001100",
    "1111110000101000",
    "1111110000010111",
    "1111110100010011",
    "1111111100011111",
    "1111111000000100",
    "1111101011011000",
    "1111011111110011",
    "1111010111011010",
    "1111010011100010",
    "1111010100101001",
    "1111011010010001",
    "1111100011011101",
    "1111101110111110",
    "1111111011011111",
    "1111111000000000",
    "1111101100011001",
    "1111100010001011",
    "1111011001101011",
    "1111010011000011",
    "1111001110010100",
    "1111001011100001",
    "1111001010100110",
    "1111001011100000",
    "1111001110000111",
    "1111010010010010",
    "1111010111110111",
    "1111011110101011",
    "1111100110100111",
    "1111101111100111",
    "1111111001110010",
    "1111111010100110",
    "1111101101010111",
    "1111011110011100",
    "1111001110010111",
    "1110111110010010",
    "1110101111110110",
    "1110100100110011",
    "1110011110011110",
    "1110011101011011",
    "1110100001010100",
    "1110101001000111",
    "1110110011100100",
    "1110111111100100",
    "1111001100101010",
    "1111011010111010",
    "1111101010101011",
    "1111111011111011",
    "1111110001111101",
    "1111100000100100",
    "1111010001101100",
    "1111000111001001",
    "1111000001111101",
    "1111000010001111",
    "1111000111001000",
    "1111001111010010",
    "1111011001011000",
    "1111100100010011",
    "1111101111010001",
    "1111111001100101",
    "1111111101100110",
    "1111110111010100",
    "1111110100011111",
    "1111110101101000",
    "1111111010100001",
    "1111111101111010",
    "1111110101100001",
    "1111101110001101",
    "1111101001110000",
    "1111101001001011",
    "1111101100110101",
    "1111110100100100",
    "1111111111111000",
    "1111110001111011",
    "1111100001111000",
    "1111010001010010",
    "1111000001110100",
    "1110110101001101",
    "1110101100111101",
    "1110101010000111",
    "1110101101000111",
    "1110110101111001",
    "1111000011110100",
    "1111010101101010",
    "1111101001101101",
    "1111111101110001",
    "1111110000010000",
    "1111100010001011",
    "1111011000110111",
    "1111010100010010",
    "1111010011100111",
    "1111010101110110",
    "1111011010000010",
    "1111011111111101",
    "1111100111101010",
    "1111110001100101",
    "1111111101110110",
    "1111110011110100",
    "1111100100011111",
    "1111010101100111",
    "1111001000101101",
    "1110111110111111",
    "1110111001000010",
    "1110110110110010",
    "1110110111100111",
    "1110111010100010",
    "1110111110101101",
    "1111000011010111",
    "1111001000000110",
    "1111001100101101",
    "1111010001001111",
    "1111010101101111",
    "1111011010001110",
    "1111011110100110",
    "1111100010101011",
    "1111100110001000",
    "1111101000110110",
    "1111101010101111",
    "1111101011111100",
    "1111101100101001",
    "1111101101001011",
    "1111101101111000",
    "1111101111001000",
    "1111110001011000",
    "1111110101001011",
    "1111111011000100",
    "1111111100011111",
    "1111110001100000",
    "1111100100011101",
    "1111010110011101",
    "1111001001010001",
    "1110111110110000",
    "1110111000100010",
    "1110110111100011",
    "1110111011110111",
    "1111000100110110",
    "1111010001010111",
    "1111100000010100",
    "1111110000101110",
    "1111111110001001",
    "1111101100111100",
    "1111011100010001",
    "1111001100111111",
    "1111000000000010",
    "1110110110010011",
    "1110110000010100",
    "1110101101111111",
    "1110101110100001",
    "1110110000100110",
    "1110110010110100",
    "1110110011111110",
    "1110110011011100",
    "1110110001001111",
    "1110101101111111",
    "1110101010101010",
    "1110101000000110",
    "1110100110111111",
    "1110100111100101",
    "1110101001101111",
    "1110101100111111",
    "1110110000111001",
    "1110110100111110",
    "1110111000110111",
    "1110111100011011",
    "1110111111101001",
    "1111000010100100",
    "1111000101001110",
    "1111000111101111",
    "1111001010000110",
    "1111001100001110",
    "1111001101111111",
    "1111001111001101",
    "1111001111101100",
    "1111001111010010",
    "1111001110000010",
    "1111001100000111",
    "1111001001111001",
    "1111000111110111",
    "1111000110101000",
    "1111000110101010",
    "1111001000010001",
    "1111001011100011",
    "1111010000001101",
    "1111010101101010",
    "1111011011001001",
    "1111011111110101",
    "1111100011000101",
    "1111100100100000",
    "1111100100010101",
    "1111100011000110",
    "1111100001110000",
    "1111100001010100",
    "1111100010110001",
    "1111100110110000",
    "1111101101011110",
    "1111110110110101",
    "1111111101100011",
    "1111110000011011",
    "1111100010101110",
    "1111010101011101",
    "1111001001101101",
    "1111000000011110",
    "1110111010010110",
    "1110110111101010",
    "1110111000010101",
    "1110111011111100",
    "1111000010000011",
    "1111001010010100",
    "1111010100100111",
    "1111100000111110",
    "1111101111010100",
    "1111111111001010",
    "1111110000011011",
    "1111100000111110",
    "1111010100000101",
    "1111001010111111",
    "1111000110011000",
    "1111000101111100",
    "1111001000101111",
    "1111001101010110",
    "1111010010011111",
    "1111010111001001",
    "1111011010111000",
    "1111011101101001",
    "1111011111110000",
    "1111100001011110",
    "1111100011001011",
    "1111100101000001",
    "1111100111001000",
    "1111101001100100",
    "1111101100011001",
    "1111101111110100",
    "1111110011111101",
    "1111111001000000",
    "1111111111000001",
    "1111111010000100",
    "1111110010100111",
    "1111101011001001",
    "1111100100001110",
    "1111011110011110",
    "1111011010001001",
    "1111010111001001",
    "1111010100111011",
    "1111010010101100",
    "1111001111100110",
    "1111001011001001",
    "1111000101010010",
    "1110111110100011",
    "1110110111111001",
    "1110110010011101",
    "1110101111001111",
    "1110101110111010",
    "1110110001100111",
    "1110110111010000",
    "1110111111011110",
    "1111001001110100",
    "1111010101101111",
    "1111100010011101",
    "1111101110110010",
    "1111111001000110",
    "1111111111101001",
    "1111111110111110",
    "1111111100010110",
    "1111110001111111",
    "1111100011010011",
    "1111010010100010",
    "1111000010010101",
    "1110110101001001",
    "1110101100110010",
    "1110101010001001",
    "1110101101001010",
    "1110110101000000",
    "1111000000010010",
    "1111001101010110",
    "1111011010100011",
    "1111100110011101",
    "1111110000001010",
    "1111110111010101",
    "1111111100001100",
    "1111111111011111",
    "1111111101110110",
    "1111111011000001",
    "1111110111100001",
    "1111110011001110",
    "1111101110010111",
    "1111101001011001",
    "1111100100110100",
    "1111100001000000",
    "1111011110010001",
    "1111011100100110",
    "1111011011111101",
    "1111011100001110",
    "1111011101001100",
    "1111011110110001",
    "1111100000111000",
    "1111100011011111",
    "1111100110100111",
    "1111101010010011",
    "1111101110101101",
    "1111110011111011",
    "1111111010000110",
    "1111111110101111",
    "1111110110101101",
    "1111101101111000",
    "1111100100011111",
    "1111011010101101",
    "1111010000110110",
    "1111000111001001",
    "1110111101110111",
    "1110110101010000",
    "1110101101011110",
    "1110100110100111",
    "1110100000101110",
    "1110011011110011",
    "1110010111111010",
    "1110010101001011",
    "1110010011110110",
    "1110010100010010",
    "1110010110111110",
    "1110011100011011",
    "1110100101001001",
    "1110110001100111",
    "1111000010000010",
    "1111010110000011",
    "1111101100100100",
    "1111111100100000",
    "1111100111111100",
    "1111011000011000",
    "1111001111100110",
    "1111001101111101",
    "1111010010001101",
    "1111011010000001",
    "1111100010110011",
    "1111101010100001",
    "1111110000010111",
    "1111110100101001",
    "1111111000011010",
    "1111111100111010",
    "1111111100111110",
    "1111110101001011",
    "1111101100010001",
    "1111100011010111",
    "1111011011101000",
    "1111010110000110",
    "1111010011010101",
    "1111010011010010",
    "1111010101011111",
    "1111011001000111",
    "1111011101001001",
    "1111100000100100",
    "1111100010101001",
    "1111100010111110",
    "1111100001100111",
    "1111011110111111",
    "1111011011101111",
    "1111011000101000",
    "1111010110011010",
    "1111010101100100",
    "1111010110011011",
    "1111011001000110",
    "1111011101010010",
    "1111100010101100",
    "1111101000110000",
    "1111101110111111",
    "1111110101000001",
    "1111111010100101",
    "1111111111100110",
    "1111111011110011",
    "1111110111100101",
    "1111110011011111",
    "1111101111011101",
    "1111101011100100",
    "1111101000000111",
    "1111100101100111",
    "1111100100101001",
    "1111100101110001",
    "1111101001010010",
    "1111101111011000",
    "1111110111111111",
    "1111111101000111",
    "1111110000011011",
    "1111100010110011",
    "1111010101011111",
    "1111001010000100",
    "1111000010001010",
    "1110111111001100",
    "1111000001111110",
    "1111001010101000",
    "1111011000011011",
    "1111101001111100",
    "1111111101001110",
    "1111110000000100",
    "1111100000001111",
    "1111010101000110",
    "1111001111110001",
    "1111010000011111",
    "1111010110101100",
    "1111100001001111",
    "1111101110011110",
    "1111111100100100",
    "1111110110010100",
    "1111101100000000",
    "1111100101101110",
    "1111100100001011",
    "1111100111011001",
    "1111101110110100",
    "1111111001010100",
    "1111111010100111",
    "1111101110101111",
    "1111100100100010",
    "1111011101001111",
    "1111011001100010",
    "1111011001100000",
    "1111011100110111",
    "1111100011000101",
    "1111101011101001",
    "1111110110000010",
    "1111111110010011",
    "1111110010001100",
    "1111100110011101",
    "1111011100000010",
    "1111010011110001",
    "1111001110001101",
    "1111001011100101",
    "1111001011110000",
    "1111001110010111",
    "1111010011000001",
    "1111011001011000",
    "1111100001010000",
    "1111101010101110",
    "1111110101111001",
    "1111111101001000",
    "1111101110101000",
    "1111011111000100",
    "1111001111011110",
    "1111000001000111",
    "1110110101010101",
    "1110101101010001",
    "1110101001011110",
    "1110101001101111",
    "1110101101001010",
    "1110110010100001",
    "1110111000101100",
    "1110111110111101",
    "1111000101011000",
    "1111001100101010",
    "1111010101110001",
    "1111100001100110",
    "1111110000011101",
    "1111111110010000",
    "1111101100011010",
    "1111011100011001",
    "1111010000100001",
    "1111001010011101",
    "1111001010100011",
    "1111010000000000",
    "1111011001010000",
    "1111100100011010",
    "1111110000000100",
    "1111111011010111",
    "1111111010000000",
    "1111110000011110",
    "1111101000100001",
    "1111100010111110",
    "1111100000101110",
    "1111100010011111",
    "1111101000010110",
    "1111110001101011",
    "1111111101000111",
    "1111110111000011",
    "1111101100100011",
    "1111100100101001",
    "1111011111110110",
    "1111011110001100",
    "1111011111001100",
    "1111100010001010",
    "1111100110011110",
    "1111101011101000",
    "1111110001011100",
    "1111110111101110",
    "1111111110011000",
    "1111111010111010",
    "1111110100110001",
    "1111101111110111",
    "1111101100111001",
    "1111101100010101",
    "1111101110010101",
    "1111110010101011",
    "1111111000101100",
    "1111111111100010",
    "1111111001101100",
    "1111110100000011",
    "1111110000010011",
    "1111101111000101",
    "1111110000110010",
    "1111110101101000",
    "1111111101100110",
    "1111110111100101",
    "1111101010100011",
    "1111011100001001",
    "1111001101100001",
    "1110111111111111",
    "1110110100101100",
    "1110101100100110",
    "1110101000001000",
    "1110100111001110",
    "1110101001100101",
    "1110101110101011",
    "1110110110001001",
    "1110111111110101",
    "1111001011101010",
    "1111011001100010",
    "1111101001000100",
    "1111111001010100",
    "1111110111000111",
    "1111101001110110",
    "1111100000010010",
    "1111011011010100",
    "1111011011001110",
    "1111011111110110",
    "1111101000110001",
    "1111110101100100",
    "1111111010011110",
    "1111101000101101",
    "1111010110111111",
    "1111000111110001",
    "1110111101010001",
    "1110111001011000",
    "1110111101000000",
    "1111001000000110",
    "1111011001100011",
    "1111101111010010",
    "1111111001101001",
    "1111100100100111",
    "1111010100101110",
    "1111001100000101",
    "1111001011100001",
    "1111010010010101",
    "1111011110100110",
    "1111101101111011",
    "1111111110001010",
    "1111110010001000",
    "1111100011101111",
    "1111010110111110",
    "1111001100000101",
    "1111000011101100",
    "1110111110101001",
    "1110111110000010",
    "1111000010011101",
    "1111001011110011",
    "1111011000111100",
    "1111100111111111",
    "1111110110110101",
    "1111111100001110",
    "1111110010010111",
    "1111101011111100",
    "1111101000110100",
    "1111101000100110",
    "1111101010110110",
    "1111101111010001",
    "1111110101101010",
    "1111111101110111",
    "1111111000010010",
    "1111101101001110",
    "1111100001011010",
    "1111010101100010",
    "1111001010010011",
    "1111000000010101",
    "1110111000001011",
    "1110110010001000",
    "1110101110010100",
    "1110101100101011",
    "1110101100111100",
    "1110101110101000",
    "1110110001010100",
    "1110110100100111",
    "1110111000010101",
    "1110111100100001",
    "1111000001011010",
    "1111000111010001",
    "1111001110011011",
    "1111010111000011",
    "1111100001010000",
    "1111101100111111",
    "1111111001101011",
    "1111111001100101",
    "1111101110001000",
    "1111100101001101",
    "1111011111110001",
    "1111011110001111",
    "1111100000001101",
    "1111100100101111",
    "1111101010011100",
    "1111110000000010",
    "1111110100011001",
    "1111110110110101",
    "1111110110111101",
    "1111110100101101",
    "1111110000010100",
    "1111101010010001",
    "1111100011010011",
    "1111011100010111",
    "1111010110011000",
    "1111010010001101",
    "1111010000010111",
    "1111010000111101",
    "1111010011110001",
    "1111011000010101",
    "1111011110001100",
    "1111100100111011",
    "1111101100011001",
    "1111110100011010",
    "1111111100110101",
    "1111111010101100",
    "1111110010110110",
    "1111101100011101",
    "1111101000011011",
    "1111100111100000",
    "1111101001111100",
    "1111101111100001",
    "1111110111011100",
    "1111111111010110",
    "1111110110001001",
    "1111101110000001",
    "1111100111110101",
    "1111100100001010",
    "1111100011010101",
    "1111100101100111",
    "1111101011001000",
    "1111110011101101",
    "1111111110111011",
    "1111110100000010",
    "1111100110011010",
    "1111011001011101",
    "1111001110010111",
    "1111000101111100",
    "1111000000011110",
    "1110111101110111",
    "1110111101100110",
    "1110111111000101",
    "1111000001101110",
    "1111000101000001",
    "1111001000101111",
    "1111001100101011",
    "1111010000110101",
    "1111010101010000",
    "1111011001111111",
    "1111011110111011",
    "1111100011111001",
    "1111101000011001",
    "1111101011110010",
    "1111101101010110",
    "1111101100011101",
    "1111101000110111",
    "1111100010111011",
    "1111011011100001",
    "1111010100000000",
    "1111001101110101",
    "1111001010010011",
    "1111001010000111",
    "1111001101011110",
    "1111010011111001",
    "1111011100100000",
    "1111100110010101",
    "1111110000101011",
    "1111111011000100",
    "1111111010110001",
    "1111110001011000",
    "1111101001100011",
    "1111100100010111",
    "1111100010111101",
    "1111100110000011",
    "1111101101101011",
    "1111111000110011",
    "1111111010001101",
    "1111101101011101",
    "1111100010110001",
    "1111011011010100",
    "1111010111101000",
    "1111010111100000",
    "1111011010010011",
    "1111011111010001",
    "1111100101101100",
    "1111101100111010",
    "1111110100011000",
    "1111111011100111",
    "1111111101110010",
    "1111111000001100",
    "1111110011100111",
    "1111101111111000",
    "1111101100101010",
    "1111101001100001",
    "1111100110000110",
    "1111100001111110",
    "1111011100111101",
    "1111010110110100",
    "1111001111100001",
    "1111000111010101",
    "1110111110101001",
    "1110110110001011",
    "1110101110101011",
    "1110101000110100",
    "1110100101000101",
    "1110100011100010",
    "1110100100000110",
    "1110100110011000",
    "1110101010000010",
    "1110101110110000",
    "1110110100010010",
    "1110111010010100",
    "1111000000011100",
    "1111000101111001",
    "1111001001110010",
    "1111001011001110",
    "1111001001100000",
    "1111000100100010",
    "1110111100101110",
    "1110110011001011",
    "1110101001010001",
    "1110100000100111",
    "1110011010100011",
    "1110011000000100",
    "1110011001101101",
    "1110011111011110",
    "1110101000110101",
    "1110110100110011",
    "1111000001110011",
    "1111001110000100",
    "1111010111110001",
    "1111011101100110",
    "1111011110111011",
    "1111011100000010",
    "1111010101110111",
    "1111001101101101",
    "1111000100101110",
    "1110111011110000",
    "1110110011010000",
    "1110101011011011",
    "1110100100011111",
    "1110011111000000",
    "1110011011110000",
    "1110011011101101",
    "1110011111100100",
    "1110100111101100",
    "1110110011101001",
    "1111000010010111",
    "1111010010011001",
    "1111100010000000",
    "1111101111101011",
    "1111111010001111",
    "1111111111000001",
    "1111111100011000",
    "1111111101101100",
    "1111111101100110",
    "1111110110010011",
    "1111101101011000",
    "1111100011110100",
    "1111011010101101",
    "1111010010111001",
    "1111001101000010",
    "1111001001100000",
    "1111001000011000",
    "1111001001100101",
    "1111001100110010",
    "1111010001100111",
    "1111010111100101",
    "1111011110000111",
    "1111100100100111",
    "1111101010100010",
    "1111101111011100",
    "1111110011001100",
    "1111110101110110",
    "1111110111101100",
    "1111111001001011",
    "1111111010100101",
    "1111111100001000",
    "1111111101110010",
    "1111111111011010",
    "1111111111001010",
    "1111111110001001",
    "1111111101011111",
    "1111111101000110",
    "1111111100101011",
    "1111111011110011",
    "1111111001111011",
    "1111110110011000",
    "1111110000100011",
    "1111101000000110",
    "1111011101001010",
    "1111010000100111",
    "1111000011111000",
    "1110111000101111",
    "1110110001000010",
    "1110101110000111",
    "1110110000101110",
    "1110111000110101",
    "1111000110000011",
    "1111010111101010",
    "1111101100111110",
    "1111111011000111",
    "1111100010010111",
    "1111001011000010",
    "1110110111100111",
    "1110101010000111",
    "1110100011100010",
    "1110100011100001",
    "1110101000010101",
    "1110101111100110",
    "1110110111000100",
    "1110111101001110",
    "1111000001011111",
    "1111000100001011",
    "1111000110000000",
    "1111000111101101",
    "1111001001111001",
    "1111001100110010",
    "1111010000011111",
    "1111010101001011",
    "1111011011000111",
    "1111100010101110",
    "1111101100011010",
    "1111111000011111",
    "1111111001000100",
    "1111101000110110",
    "1111010111110010",
    "1111000111010011",
    "1110111000110010",
    "1110101101100001",
    "1110100110001110",
    "1110100010111101",
    "1110100011001111",
    "1110100110001011",
    "1110101010110101",
    "1110110000100001",
    "1110110110101101",
    "1110111101000010",
    "1111000011001111",
    "1111001000111111",
    "1111001110000010",
    "1111010010000010",
    "1111010100110100",
    "1111010110011111",
    "1111010111011000",
    "1111011000001000",
    "1111011001100011",
    "1111011100100000",
    "1111100001011100",
    "1111101000011101",
    "1111110001001000",
    "1111111010100100",
    "1111111100010000",
    "1111110100100001",
    "1111101110111100",
    "1111101011111011",
    "1111101011011111",
    "1111101101011100",
    "1111110001100101",
    "1111110111110101",
    "1111111111101110",
    "1111110101001010",
    "1111101000101001",
    "1111011010111010",
    "1111001101001111",
    "1111000001010100",
    "1110111000111111",
    "1110110101110110",
    "1110111000101111",
    "1111000001100111",
    "1111001111010111",
    "1111100000000000",
    "1111110001010101",
    "1111111110101011",
    "1111110001100010",
    "1111100111110101",
    "1111100001011010",
    "1111011101101110",
    "1111011100000010",
    "1111011011110010",
    "1111011100101101",
    "1111011110111010",
    "1111100010101001",
    "1111101000000100",
    "1111101111001000",
    "1111110111100010",
    "1111111111010001",
    "1111110110000001",
    "1111101101010001",
    "1111100101100000",
    "1111011110111011",
    "1111011001011110",
    "1111010100110011",
    "1111010000011001",
    "1111001011110000",
    "1111000110011101",
    "1111000000001100",
    "1110111000111100",
    "1110110000110101",
    "1110101000001000",
    "1110011111000101",
    "1110010101111011",
    "1110001100110011",
    "1110000011111100",
    "1101111011100011",
    "1101110011111110",
    "1101101101101000",
    "1101101001000100",
    "1101100110101111",
    "1101100111000011",
    "1101101010000111",
    "1101101111110011",
    "1101110111101100",
    "1110000001001101",
    "1110001011110111",
    "1110010111010011",
    "1110100011101001",
    "1110110001001100",
    "1111000000010001",
    "1111010000110011",
    "1111100010000011",
    "1111110010100110",
    "1111111111010101",
    "1111110101101000",
    "1111110001100011",
    "1111110011100100",
    "1111111011000110",
    "1111111001001011",
    "1111101011001111",
    "1111011101001110",
    "1111010001010100",
    "1111001001010001",
    "1111000110011101",
    "1111001001010101",
    "1111010001011111",
    "1111011101101011",
    "1111101011111010",
    "1111111001110110",
    "1111111010100001",
    "1111110010101110",
    "1111101111010110",
    "1111110000000101",
    "1111110100000110",
    "1111111010010110",
    "1111111110001110",
    "1111110110101001",
    "1111101111110100",
    "1111101010011110",
    "1111100111010000",
    "1111100110011101",
    "1111100111111011",
    "1111101011000010",
    "1111101110110111",
    "1111110010011000",
    "1111110100110100",
    "1111110101111101",
    "1111110110000010",
    "1111110101101110",
    "1111110101110010",
    "1111110110110001",
    "1111111000111000",
    "1111111011110111",
    "1111111111001000",
    "1111111110000011",
    "1111111100011111",
    "1111111100110110",
    "1111111111100111",
    "1111111010111110",
    "1111110011000011",
    "1111101001001000",
    "1111011110000100",
    "1111010010111101",
    "1111001001000001",
    "1111000001010000",
    "1110111100010110",
    "1110111010011110",
    "1110111011011110",
    "1110111110111011",
    "1111000100100010",
    "1111001100000100",
    "1111010101101010",
    "1111100001110011",
    "1111110001000001",
    "1111111011111110",
    "1111100101001000",
    "1111001011001100",
    "1110110000010010",
    "1110010111010011",
    "1110000011001011",
    "1101110110000011",
    "1101110000100111",
    "1101110010000110",
    "1101111000100101",
    "1110000001111110",
    "1110001100101110",
    "1110011000010001",
    "1110100100101110",
    "1110110010001111",
    "1111000000011110",
    "1111001110010110",
    "1111011010001011",
    "1111100010001111",
    "1111100101011011",
    "1111100011110011",
    "1111011110010111",
    "1111010110111111",
    "1111001111101100",
    "1111001010001001",
    "1111000111010110",
    "1111000111111001",
    "1111001011110101",
    "1111010010111110",
    "1111011100110010",
    "1111101000011011",
    "1111110100101101",
    "1111111111101100",
    "1111110110001010",
    "1111101111101001",
    "1111101100101011",
    "1111101101001110",
    "1111110000110101",
    "1111110110110111",
    "1111111110110010",
    "1111110111110011",
    "1111101101010000",
    "1111100001111001",
    "1111010110010110",
    "1111001011011001",
    "1111000010000011",
    "1110111011010001",
    "1110110111101101",
    "1110110111110100",
    "1110111011100101",
    "1111000010101111",
    "1111001100110111",
    "1111011001010000",
    "1111100111000010",
    "1111110101001010",
    "1111111101011000",
    "1111110001100111",
    "1111101000001111",
    "1111100001100110",
    "1111011101110010",
    "1111011100100011",
    "1111011101100100",
    "1111100000100100",
    "1111100101010111",
    "1111101011110100",
    "1111110011111001",
    "1111111101100011",
    "1111110111001110",
    "1111101010101111",
    "1111011101100011",
    "1111010000100110",
    "1111000101000101",
    "1110111100001010",
    "1110110110110010",
    "1110110101011010",
    "1110110111111100",
    "1110111101101011",
    "1111000101100100",
    "1111001110001111",
    "1111010110001101",
    "1111011011111000",
    "1111011101110101",
    "1111011011000001",
    "1111010011000001",
    "1111000110100111",
    "1110110111011111",
    "1110101000001001",
    "1110011011001110",
    "1110010010111011",
    "1110010000011100",
    "1110010011111110",
    "1110011100110111",
    "1110101010000111",
    "1110111010110111",
    "1111001110011111",
    "1111100100011000",
    "1111111011011101",
    "1111101101111011",
    "1111011010000100",
    "1111001011000110",
    "1111000010011100",
    "1111000000011001",
    "1111000011110110",
    "1111001010111010",
    "1111010011011010",
    "1111011011101111",
    "1111100011001011",
    "1111101001111011",
    "1111110000101011",
    "1111111000001000",
    "1111111111010001",
    "1111110101101011",
    "1111101011100000",
    "1111100001011110",
    "1111011000010110",
    "1111010000111000",
    "1111001011101010",
    "1111001001000111",
    "1111001001011011",
    "1111001100011110",
    "1111010001110100",
    "1111011000110101",
    "1111100000111000",
    "1111101001100011",
    "1111110010101010",
    "1111111100001101",
    "1111111001110110",
    "1111101111111001",
    "1111100110011011",
    "1111011110001100",
    "1111010111111010",
    "1111010100000001",
    "1111010010100111",
    "1111010011010111",
    "1111010101101111",
    "1111011001001110",
    "1111011101010110",
    "1111100001110000",
    "1111100110001000",
    "1111101010000001",
    "1111101100110101",
    "1111101101111111",
    "1111101100111110",
    "1111101001101110",
    "1111100100101010",
    "1111011110101110",
    "1111011001001001",
    "1111010101000110",
    "1111010011011111",
    "1111010100110001",
    "1111011000111001",
    "1111011111011111",
    "1111100111111111",
    "1111110001110010",
    "1111111100011001",
    "1111111000100011",
    "1111101101100011",
    "1111100011000101",
    "1111011001110000",
    "1111010010010111",
    "1111001101101001",
    "1111001100001001",
    "1111001110000010",
    "1111010011000011",
    "1111011010011011",
    "1111100011001101",
    "1111101100010111",
    "1111110100111111",
    "1111111100011111",
    "1111111101011111",
    "1111111001001100",
    "1111110110100100",
    "1111110101100110",
    "1111110110001011",
    "1111111000000001",
    "1111111010110011",
    "1111111101111010",
    "1111111111001110",
    "1111111101010001",
    "1111111100100000",
    "1111111101000000",
    "1111111110011110",
    "1111111111100000",
    "1111111101011010",
    "1111111011100001",
    "1111111001111100",
    "1111111000100101",
    "1111110111010101",
    "1111110110000001",
    "1111110100101011",
    "1111110011011001",
    "1111110010010010",
    "1111110001100001",
    "1111110001001010",
    "1111110001010000",
    "1111110001110100",
    "1111110010110110",
    "1111110100010101",
    "1111110110010101",
    "1111111000111010",
    "1111111100000011",
    "1111111111101110",
    "1111111100001110",
    "1111111000010011",
    "1111110101000110",
    "1111110011010100",
    "1111110011110001",
    "1111110111000010",
    "1111111101001110",
    "1111111010000110",
    "1111110000000110",
    "1111100110010010",
    "1111011110010111",
    "1111011001110101",
    "1111011001101010",
    "1111011110001101",
    "1111100111100001",
    "1111110101010010",
    "1111111000111111",
    "1111100100011111",
    "1111001111000010",
    "1110111010111101",
    "1110101010101011",
    "1110100000000000",
    "1110011011101000",
    "1110011101000100",
    "1110100010101110",
    "1110101010100101",
    "1110110010111001",
    "1110111010101011",
    "1111000001100111",
    "1111000111111010",
    "1111001101111010",
    "1111010011110100",
    "1111011001100111",
    "1111011111000010",
    "1111100011111100",
    "1111101000010110",
    "1111101100100001",
    "1111110000111010",
    "1111110110000001",
    "1111111100010000",
    "1111111100000111",
    "1111110011000110",
    "1111101000110111",
    "1111011101111011",
    "1111010011001000",
    "1111001001011000",
    "1111000001100001",
    "1110111011111100",
    "1110111000101000",
    "1110110111001001",
    "1110110110110100",
    "1110110111000110",
    "1110110111101010",
    "1110111000011011",
    "1110111001100011",
    "1110111011001110",
    "1110111101100000",
    "1111000000010010",
    "1111000011010111",
    "1111000110010110",
    "1111001001001011",
    "1111001011110101",
    "1111001110101101",
    "1111010010010111",
    "1111010111011011",
    "1111011110011100",
    "1111100111101011",
    "1111110011000101",
    "1111111111111100",
    "1111110010101011",
    "1111100110100101",
    "1111011101001010",
    "1111010111011101",
    "1111010101110001",
    "1111010111100011",
    "1111011011110000",
    "1111100001000000",
    "1111100110001000",
    "1111101010011001",
    "1111101101100011",
    "1111101111101100",
    "1111110001000101",
    "1111110001111000",
    "1111110010000111",
    "1111110001101011",
    "1111110000011101",
    "1111101110011100",
    "1111101011110000",
    "1111101000101010",
    "1111100101011111",
    "1111100010100010",
    "1111100000001010",
    "1111011110100110",
    "1111011110001101",
    "1111011111010100",
    "1111100010000011",
    "1111100110011111",
    "1111101100011001",
    "1111110011011100",
    "1111111011001000",
    "1111111100111111",
    "1111110101011101",
    "1111101110100101",
    "1111101000100100",
    "1111100011100010",
    "1111011111100001",
    "1111011100011011",
    "1111011010000111",
    "1111011000010001",
    "1111010110100101",
    "1111010100110001",
    "1111010010101011",
    "1111010000010101",
    "1111001110000111",
    "1111001100011011",
    "1111001011101010",
    "1111001100000100",
    "1111001101101101",
    "1111010000011010",
    "1111010011111000",
    "1111010111110010",
    "1111011011110101",
    "1111011111110001",
    "1111100011011111",
    "1111100110111001",
    "1111101001111101",
    "1111101100110011",
    "1111101111100010",
    "1111110010011010",
    "1111110101110100",
    "1111111010000011",
    "1111111111010101",
    "1111111010011000",
    "1111110011011111",
    "1111101100101001",
    "1111100110101010",
    "1111100010011010",
    "1111100000011111",
    "1111100001010100",
    "1111100100111001",
    "1111101011001010",
    "1111110100000000",
    "1111111111010011",
    "1111110011000001",
    "1111100011100100",
    "1111010011011010",
    "1111000100010000",
    "1110111000000011",
    "1110110000011100",
    "1110101110001101",
    "1110110001000010",
    "1110110111100011",
    "1110111111110110",
    "1111000111111111",
    "1111001110100100",
    "1111010010111000",
    "1111010100110011",
    "1111010100101010",
    "1111010011000001",
    "1111010000011001",
    "1111001101010110",
    "1111001010011011",
    "1111001000010000",
    "1111000111010101",
    "1111001000001000",
    "1111001010101101",
    "1111001110110101",
    "1111010011111011",
    "1111011001000100",
    "1111011101011110",
    "1111100000010111",
    "1111100001010000",
    "1111100000000010",
    "1111011100110011",
    "1111011000000100",
    "1111010010100010",
    "1111001100111111",
    "1111001000001011",
    "1111000100101001",
    "1111000010101100",
    "1111000010010111",
    "1111000011010011",
    "1111000101001001",
    "1111000111011010",
    "1111001001101111",
    "1111001011111101",
    "1111001110000000",
    "1111001111111010",
    "1111010001100110",
    "1111010011000011",
    "1111010100000011",
    "1111010100100010",
    "1111010100100000",
    "1111010100010010",
    "1111010100010010",
    "1111010101001000",
    "1111010111011000",
    "1111011011100110",
    "1111100010001010",
    "1111101011010101",
    "1111110111001011",
    "1111111010101000",
    "1111101010111110",
    "1111011011000010",
    "1111001100011001",
    "1111000000100111",
    "1110111001000001",
    "1110110110010101",
    "1110111000111100",
    "1111000000110001",
    "1111001101100100",
    "1111011110100110",
    "1111110010011011",
    "1111111001001000",
    "1111100110110000",
    "1111011000110010",
    "1111010000110001",
    "1111001110110011",
    "1111010001100111",
    "1111010111000110",
    "1111011101000010",
    "1111100001111000",
    "1111100101000110",
    "1111100111000101",
    "1111101000101101",
    "1111101010110000",
    "1111101101101010",
    "1111110001001100",
    "1111110100101111",
    "1111110111100100",
    "1111111001001001",
    "1111111001001100",
    "1111110111110110",
    "1111110101010110",
    "1111110010000000",
    "1111101110010001",
    "1111101010100110",
    "1111100111101000",
    "1111100101111110",
    "1111100110001001",
    "1111101000011110",
    "1111101100111011",
    "1111110011001110",
    "1111111010110111",
    "1111111100110010",
    "1111110100011100",
    "1111101100101000",
    "1111100101101110",
    "1111011111111011",
    "1111011011010100",
    "1111010111110111",
    "1111010101100101",
    "1111010100011010",
    "1111010100010011",
    "1111010101001101",
    "1111010110111111",
    "1111011001100011",
    "1111011100110010",
    "1111100000010111",
    "1111100011110011",
    "1111100110011110",
    "1111100111101001",
    "1111100110101000",
    "1111100010111110",
    "1111011100011110",
    "1111010011001011",
    "1111000111100000",
    "1110111010000110",
    "1110101011111100",
    "1110011110010100",
    "1110010010101110",
    "1110001010100110",
    "1110000111001001",
    "1110001001010000",
    "1110010001000010",
    "1110011101111111",
    "1110101110101000",
    "1111000000110101",
    "1111010010000010",
    "1111011111101110",
    "1111101000000101",
    "1111101010010011",
    "1111100110101001",
    "1111011110001100",
    "1111010010010100",
    "1111000100100101",
    "1110110110011000",
    "1110101001000001",
    "1110011101110000",
    "1110010101101010",
    "1110010001100001",
    "1110010001101100",
    "1110010101110111",
    "1110011101001001",
    "1110100110000100",
    "1110101111001000",
    "1110110110111011",
    "1110111100011110",
    "1110111111011001",
    "1110111111101110",
    "1110111101111111",
    "1110111010110010",
    "1110110110101111",
    "1110110010011010",
    "1110101110001010",
    "1110101010010100",
    "1110100111000100",
    "1110100100011101",
    "1110100010100110",
    "1110100001100010",
    "1110100001011110",
    "1110100010100100",
    "1110100101000101",
    "1110101001001011",
    "1110101110111000",
    "1110110110001110",
    "1110111111000010",
    "1111001001001011",
    "1111010100010111",
    "1111100000010001",
    "1111101100011111",
    "1111111000100110",
    "1111111011110110",
    "1111110001011101",
    "1111101000101010",
    "1111100001110011",
    "1111011101000101",
    "1111011010100011",
    "1111011010000010",
    "1111011011011000",
    "1111011110011001",
    "1111100011000011",
    "1111101001011101",
    "1111110001111001",
    "1111111100100111",
    "1111110110011100",
    "1111100111111110",
    "1111011001001100",
    "1111001011101111",
    "1111000001001111",
    "1110111010111000",
    "1110111001000111",
    "1110111011101011",
    "1111000001110011",
    "1111001010100010",
    "1111010101001000",
    "1111100000111011",
    "1111101101011000",
    "1111111001100111",
    "1111111011010111",
    "1111110010110100",
    "1111101101101101",
    "1111101100100100",
    "1111101111010001",
    "1111110101000101",
    "1111111100110100",
    "1111111010110110",
    "1111110011001001",
    "1111101100111001",
    "1111101000100101",
    "1111100110010110",
    "1111100110001001",
    "1111100111110000",
    "1111101010101111",
    "1111101110101011",
    "1111110011000100",
    "1111110111011100",
    "1111111011010101",
    "1111111110010111",
    "1111111111110000",
    "1111111111010001",
    "1111111111101001",
    "1111111101000100",
    "1111111001000011",
    "1111110011110110",
    "1111101101110101",
    "1111100111100001",
    "1111100001100001",
    "1111011100011110",
    "1111011000111111",
    "1111010111100101",
    "1111011000110000",
    "1111011100111101",
    "1111100100011010",
    "1111101111001100",
    "1111111101000111",
    "1111110010010000",
    "1111011111111000",
    "1111001100111000",
    "1110111010101010",
    "1110101010011110",
    "1110011101010110",
    "1110010011110100",
    "1110001101111011",
    "1110001011010001",
    "1110001011001100",
    "1110001101000010",
    "1110010000010101",
    "1110010100111100",
    "1110011011000001",
    "1110100010101111",
    "1110101100010111",
    "1110110111110010",
    "1111000100011111",
    "1111010001011001",
    "1111011101001010",
    "1111100110011011",
    "1111101100000111",
    "1111101101101110",
    "1111101011100100",
    "1111100110101001",
    "1111100000101011",
    "1111011011110010",
    "1111011001111111",
    "1111011100111101",
    "1111100101011010",
    "1111110010110001",
    "1111111100101001",
    "1111101011011111",
    "1111011100011100",
    "1111010001101100",
    "1111001100010100",
    "1111001100001111",
    "1111010000010101",
    "1111010111001011",
    "1111011111010001",
    "1111100111110000",
    "1111110000010101",
    "1111111001001010",
    "1111111101100000",
    "1111110011101011",
    "1111101001101100",
    "1111100000010010",
    "1111011000001100",
    "1111010010000101",
    "1111001110000101",
    "1111001011111111",
    "1111001011001110",
    "1111001011001110",
    "1111001011011110",
    "1111001011110101",
    "1111001100010111",
    "1111001101011100",
    "1111001111010010",
    "1111010010000110",
    "1111010101110110",
    "1111011010001100",
    "1111011110101001",
    "1111100010101111",
    "1111100101111110",
    "1111101000000001",
    "1111101000101111",
    "1111101000001000",
    "1111100110010000",
    "1111100011011000",
    "1111011111101110",
    "1111011011100000",
    "1111010110111100",
    "1111010010001000",
    "1111001101001001",
    "1111001000000011",
    "1111000011000001",
    "1110111110010110",
    "1110111010011011",
    "1110110111110101",
    "1110110111001101",
    "1110111000111111",
    "1110111101100110",
    "1111000100111110",
    "1111001110101001",
    "1111011001101000",
    "1111100100101001",
    "1111101110010010",
    "1111110101010001",
    "1111111000110010",
    "1111111000100111",
    "1111110100111111",
    "1111101110100110",
    "1111100110010011",
    "1111011101001111",
    "1111010100011111",
    "1111001101000101",
    "1111000111111110",
    "1111000101101111",
    "1111000110101000",
    "1111001010011011",
    "1111010000100110",
    "1111011000010110",
    "1111100000110011",
    "1111101001000101",
    "1111110000011011",
    "1111110110000101",
    "1111111001011001",
    "1111111001110010",
    "1111110110110101",
    "1111110000010101",
    "1111100110100001",
    "1111011010000010",
    "1111001100000010",
    "1110111101110010",
    "1110110000101001",
    "1110100101101111",
    "1110011101110011",
    "1110011001001100",
    "1110010111111110",
    "1110011001111101",
    "1110011110111011",
    "1110100110100000",
    "1110110000001010",
    "1110111011001100",
    "1111000110101100",
    "1111010001110000",
    "1111011011100001",
    "1111100011011111",
    "1111101001010110",
    "1111101101001111",
    "1111101111011011",
    "1111110000011001",
    "1111110000100101",
    "1111110000011101",
    "1111110000011111",
    "1111110001001011",
    "1111110010111100",
    "1111110110001001",
    "1111111010111001",
    "1111111110111011",
    "1111110111110110",
    "1111110000011100",
    "1111101001010111",
    "1111100011001011",
    "1111011110001100",
    "1111011010100101",
    "1111011000001110",
    "1111010111000001",
    "1111010110110010",
    "1111010111100011",
    "1111011001011011",
    "1111011100101011",
    "1111100001110001",
    "1111101001000110",
    "1111110010110011",
    "1111111110011111",
    "1111110100110000",
    "1111101000100001",
    "1111011110011111",
    "1111011000001100",
    "1111010110101100",
    "1111011010001100",
    "1111100010011001",
    "1111101110100111",
    "1111111110010011",
    "1111101110111111",
    "1111011001111101",
    "1111000011111000",
    "1110101110100011",
    "1110011100010111",
    "1110001111011010",
    "1110001001000100",
    "1110001001010110",
    "1110001111000010",
    "1110010111111111",
    "1110100001111101",
    "1110101011000010",
    "1110110010010000",
    "1110110111010001",
    "1110111010010011",
    "1110111011110011",
    "1110111100010100",
    "1110111100010110",
    "1110111100010100",
    "1110111100110011",
    "1110111110010111",
    "1111000001100110",
    "1111000110111001",
    "1111001110100001",
    "1111011000010000",
    "1111100011100110",
    "1111101111101111",
    "1111111011101100",
    "1111111001100111",
    "1111110001001100",
    "1111101011101000",
    "1111101001001001",
    "1111101001011001",
    "1111101011101111",
    "1111101111011010",
    "1111110011110000",
    "1111111000010010",
    "1111111100111000",
    "1111111110011110",
    "1111111001111000",
    "1111110101100001",
    "1111110001110100",
    "1111101111010110",
    "1111101110100101",
    "1111101111110011",
    "1111110010111000",
    "1111110111010100",
    "1111111100010011",
    "1111111110111110",
    "1111111011010001",
    "1111111000111111",
    "1111111000001110",
    "1111111000110110",
    "1111111010100011",
    "1111111100110111",
    "1111111111001110",
    "1111111111000011",
    "1111111110110100",
    "1111111111001111",
    "1111111010110000",
    "1111110011101010",
    "1111101010100100",
    "1111100000100100",
    "1111010111000100",
    "1111001111011100",
    "1111001010101010",
    "1111001001001100",
    "1111001010111000",
    "1111001111001101",
    "1111010101100010",
    "1111011101010001",
    "1111100110001000",
    "1111110000000000",
    "1111111011000001",
    "1111111000110011",
    "1111101011101100",
    "1111011110000101",
    "1111010000110011",
    "1111000100110100",
    "1110111011000111",
    "1110110100011101",
    "1110110001000011",
    "1110110000101110",
    "1110110010110100",
    "1110110110100010",
    "1110111011000110",
    "1110111111111011",
    "1111000100101111",
    "1111001001100000",
    "1111001110010001",
    "1111010011001010",
    "1111011000001110",
    "1111011101100011",
    "1111100011001111",
    "1111101001010110",
    "1111101111111011",
    "1111110110111011",
    "1111111110001000",
    "1111111010110000",
    "1111110100010000",
    "1111101110110010",
    "1111101010101111",
    "1111101000010001",
    "1111100111010010",
    "1111100111100100",
    "1111101000110000",
    "1111101010011101",
    "1111101100011001",
    "1111101110011101",
    "1111110000101001",
    "1111110011000111",
    "1111110101111111",
    "1111111001011110",
    "1111111101101110",
    "1111111101000011",
    "1111110110110001",
    "1111101111001110",
    "1111100110011000",
    "1111011100010111",
    "1111010001101110",
    "1111000111010110",
    "1110111110100011",
    "1110111000101100",
    "1110110110111111",
    "1110111010010001",
    "1111000010100100",
    "1111001111001100",
    "1111011110101000",
    "1111101110110100",
    "1111111101101101",
    "1111110110011110",
    "1111101110110011",
    "1111101011011101",
    "1111101011110100",
    "1111101110110001",
    "1111110011000101",
    "1111110111101110",
    "1111111100000011",
    "1111111111101110",
    "1111111101010000",
    "1111111010111001",
    "1111111000111110",
    "1111110111001110",
    "1111110101010010",
    "1111110010101011",
    "1111101110110101",
    "1111101001010101",
    "1111100001111011",
    "1111011000110101",
    "1111001110110000",
    "1111000100100111",
    "1110111011100000",
    "1110110100010010",
    "1110101111100011",
    "1110101101011011",
    "1110101101101101",
    "1110110000000000",
    "1110110011111000",
    "1110111000111110",
    "1110111111000100",
    "1111000110000100",
    "1111001101111000",
    "1111010110010110",
    "1111011111010010",
    "1111101000011111",
    "1111110001110100",
    "1111111011010001",
    "1111111010111111",
    "1111110000111000",
    "1111100110011000",
    "1111011011101010",
    "1111010001001010",
    "1111000111011011",
    "1110111111000000",
    "1110111000010011",
    "1110110011010111",
    "1110110000001010",
    "1110101110011011",
    "1110101101111101",
    "1110101110101001",
    "1110110000100100",
    "1110110011111110",
    "1110111001001011",
    "1111000000100110",
    "1111001010101000",
    "1111010111100101",
    "1111100111100011",
    "1111111010001010",
    "1111110001011111",
    "1111011100111111",
    "1111001010010110",
    "1110111011101010",
    "1110110010100110",
    "1110101111111011",
    "1110110011010111",
    "1110111011101010",
    "1111000111000100",
    "1111010011101110",
    "1111100000000101",
    "1111101011000001",
    "1111110011110100",
    "1111111001111101",
    "1111111101000100",
    "1111111100110101",
    "1111111001010110",
    "1111110011000100",
    "1111101010111001",
    "1111100010000000",
    "1111011001100101",
    "1111010010100010",
    "1111001101011100",
    "1111001010011000",
    "1111001001001100",
    "1111001001101010",
    "1111001011100011",
    "1111001110110001",
    "1111010011001010",
    "1111011000010011",
    "1111011101101001",
    "1111100010011101",
    "1111100110000000",
    "1111100111101000",
    "1111100111001011",
    "1111100100110001",
    "1111100000111001",
    "1111011100001110",
    "1111010111011000",
    "1111010011000011",
    "1111001111101110",
    "1111001101110101",
    "1111001101110010",
    "1111001111110101",
    "1111010100001000",
    "1111011010101011",
    "1111100011010011",
    "1111101101101010",
    "1111111001001110",
    "1111111010011101",
    "1111101101111110",
    "1111100001100110",
    "1111010101100010",
    "1111001001111001",
    "1110111110110101",
    "1110110100101010",
    "1110101011111100",
    "1110100101010101",
    "1110100001011110",
    "1110100000110110",
    "1110100011100111",
    "1110101001101011",
    "1110110010101111",
    "1110111110011100",
    "1111001100001111",
    "1111011011100000",
    "1111101011001101",
    "1111111010000110",
    "1111111001001101",
    "1111110000000010",
    "1111101011001000",
    "1111101010100010",
    "1111101101100111",
    "1111110011001010",
    "1111111001101001",
    "1111111111011010",
    "1111111100110101",
    "1111111100001010",
    "1111111110111000",
    "1111111011010010",
    "1111110011010101",
    "1111101010110000",
    "1111100011001011",
    "1111011110000100",
    "1111011100010111",
    "1111011110010111",
    "1111100011100110",
    "1111101011010000",
    "1111110100010111",
    "1111111110000110",
    "1111111000000110",
    "1111101110101000",
    "1111100101100111",
    "1111011101001010",
    "1111010101011000",
    "1111001110010111",
    "1111001000001110",
    "1111000010111011",
    "1110111110011110",
    "1110111010110010",
    "1110110111110111",
    "1110110101101010",
    "1110110100010011",
    "1110110011110100",
    "1110110100010011",
    "1110110101110100",
    "1110111000010001",
    "1110111011100101",
    "1110111111011110",
    "1111000011101010",
    "1111000111111001",
    "1111001011101011",
    "1111001110101000",
    "1111010000001111",
    "1111010000000111",
    "1111001101111000",
    "1111001001011101",
    "1111000010111110",
    "1110111010111101",
    "1110110010000000",
    "1110101000111100",
    "1110100000100100",
    "1110011001100101",
    "1110010100100100",
    "1110010001111011",
    "1110010010000010",
    "1110010101001011",
    "1110011011101111",
    "1110100110000000",
    "1110110100000101",
    "1111000101100101",
    "1111011001011101",
    "1111101101111111",
    "1111111110110110",
    "1111101110111010",
    "1111100011010011",
    "1111011100001110",
    "1111011000110111",
    "1111010111111110",
    "1111011000010001",
    "1111011000111010",
    "1111011001101011",
    "1111011010111010",
    "1111011101000101",
    "1111100000100100",
    "1111100101010010",
    "1111101010100011",
    "1111101111011110",
    "1111110011000100",
    "1111110100101001",
    "1111110100000010",
    "1111110001100111",
    "1111101110001100",
    "1111101010110111",
    "1111101000110000",
    "1111101000110111",
    "1111101011111110",
    "1111110010100100",
    "1111111100101100",
    "1111110110000011",
    "1111100110101011",
    "1111010110011101",
    "1111000110111011",
    "1110111001011011",
    "1110101111000101",
    "1110101000011101",
    "1110100101100010",
    "1110100110000011",
    "1110101001011101",
    "1110101111000111",
    "1110110110100000",
    "1110111111000100",
    "1111001000010101",
    "1111010001110110",
    "1111011011001110",
    "1111100100000011",
    "1111101100000110",
    "1111110011001001",
    "1111111001000110",
    "1111111110000010",
    "1111111101111010",
    "1111111010101100",
    "1111111000001010",
    "1111110110010001",
    "1111110100111011",
    "1111110100000100",
    "1111110011100111",
    "1111110011011101",
    "1111110011011110",
    "1111110011100110",
    "1111110011101111",
    "1111110011110100",
    "1111110011110010",
    "1111110011100000",
    "1111110010110110",
    "1111110001101100",
    "1111110000000100",
    "1111101110001000",
    "1111101100001111",
    "1111101010111101",
    "1111101010111000",
    "1111101100101101",
    "1111110001000111",
    "1111111000100111",
    "1111111100101010",
    "1111101111100011",
    "1111100001100100",
    "1111010100110001",
    "1111001011010100",
    "1111000110101000",
    "1111000111010011",
    "1111001100101101",
    "1111010101101001",
    "1111100000101110",
    "1111101101000001",
    "1111111010001011",
    "1111110111110111",
    "1111101001100001",
    "1111011011101011",
    "1111001111111000",
    "1111000111111110",
    "1111000101011111",
    "1111001001000100",
    "1111010010010101",
    "1111011111110000",
    "1111101111001110",
    "1111111110100010",
    "1111110100000100",
    "1111101001101111",
    "1111100010110011",
    "1111011110111111",
    "1111011101101101",
    "1111011110000111",
    "1111011111010111",
    "1111100000110110",
    "1111100010001101",
    "1111100011010101",
    "1111100100010101",
    "1111100101011010",
    "1111100110101101",
    "1111101000010000",
    "1111101001110101",
    "1111101011001001",
    "1111101011110110",
    "1111101011101011",
    "1111101010100011",
    "1111101000100101",
    "1111100110000000",
    "1111100011000101",
    "1111100000001000",
    "1111011101010111",
    "1111011011000010",
    "1111011001011000",
    "1111011000100101",
    "1111011000111001",
    "1111011010010110",
    "1111011100111111",
    "1111100000100011",
    "1111100100110100",
    "1111101001100010",
    "1111101110101000",
    "1111110100000100",
    "1111111001111111",
    "1111111111011011",
    "1111111000000110",
    "1111101111111011",
    "1111100110111011",
    "1111011101010111",
    "1111010011110100",
    "1111001011000010",
    "1111000011111000",
    "1110111111000100",
    "1110111100111111",
    "1110111101101000",
    "1111000000011100",
    "1111000100101100",
    "1111001001011101",
    "1111001101110011",
    "1111010000111101",
    "1111010010010100",
    "1111010001011110",
    "1111001110010110",
    "1111001001000111",
    "1111000010001111",
    "1110111010010011",
    "1110110010000011",
    "1110101010000111",
    "1110100010111011",
    "1110011100110010",
    "1110010111111001",
    "1110010100011010",
    "1110010010011100",
    "1110010010000101",
    "1110010011011100",
    "1110010110010011",
    "1110011010010110",
    "1110011110111101",
    "1110100011100001",
    "1110100111011011",
    "1110101010010001",
    "1110101011111111",
    "1110101100101101",
    "1110101100110101",
    "1110101100111010",
    "1110101101010111",
    "1110101110101000",
    "1110110000111011",
    "1110110100100000",
    "1110111001100000",
    "1111000000000000",
    "1111000111111110",
    "1111010001000111",
    "1111011010110000",
    "1111100100000110",
    "1111101100001011",
    "1111110010001010",
    "1111110101101011",
    "1111110110101101",
    "1111110101101110",
    "1111110011011100",
    "1111110000100111",
    "1111101101111101",
    "1111101011111000",
    "1111101010101010",
    "1111101010010011",
    "1111101010101111",
    "1111101011101011",
    "1111101100110001",
    "1111101101100101",
    "1111101101110001",
    "1111101101000110",
    "1111101011100100",
    "1111101001011111",
    "1111100111100010",
    "1111100110100001",
    "1111100111010111",
    "1111101010110000",
    "1111110000111101",
    "1111111001101001",
    "1111111100000100",
    "1111110001101010",
    "1111101000100101",
    "1111100010000101",
    "1111011110111101",
    "1111011111010111",
    "1111100011000011",
    "1111101001100101",
    "1111110010011100",
    "1111111101001111",
    "1111110110011001",
    "1111101001001101",
    "1111011100001110",
    "1111010000110101",
    "1111001000011000",
    "1111000011111001",
    "1111000011100100",
    "1111000110101100",
    "1111001011111010",
    "1111010001100010",
    "1111010110001000",
    "1111011000110111",
    "1111011001101010",
    "1111011001000001",
    "1111010111101111",
    "1111010110100101",
    "1111010110001001",
    "1111010110110100",
    "1111011000101111",
    "1111011100000001",
    "1111100000110011",
    "1111100111010000",
    "1111101111100011",
    "1111111001101001",
    "1111111010110101",
    "1111101110101101",
    "1111100010111101",
    "1111011000101000",
    "1111010000101001",
    "1111001011011011",
    "1111001001000001",
    "1111001000111111",
    "1111001010110000",
    "1111001101101000",
    "1111010001000111",
    "1111010100111011",
    "1111011001000010",
    "1111011101100000",
    "1111100010010000",
    "1111100111001101",
    "1111101011111110",
    "1111110000001000",
    "1111110011001001",
    "1111110100101111",
    "1111110100111011",
    "1111110100001000",
    "1111110011000011",
    "1111110010100100",
    "1111110011011110",
    "1111110110010001",
    "1111111011001000",
    "1111111110001100",
    "1111110110011000",
    "1111101110011000",
    "1111100111001101",
    "1111100001110001",
    "1111011110110001",
    "1111011110011100",
    "1111100000100100",
    "1111100100101110",
    "1111101010001001",
    "1111110000001010",
    "1111110110000111",
    "1111111011011101",
    "1111111111110010",
    "1111111101001011",
    "1111111011110000",
    "1111111100000000",
    "1111111101111010",
    "1111111110101011",
    "1111111010001011",
    "1111110100111110",
    "1111101111100010",
    "1111101010001110",
    "1111100101011000",
    "1111100001010100",
    "1111011110001100",
    "1111011100001111",
    "1111011011101011",
    "1111011100101010",
    "1111011111001100",
    "1111100011001011",
    "1111101000011111",
    "1111101110101111",
    "1111110101100000",
    "1111111100010110",
    "1111111101000100",
    "1111110111000101",
    "1111110001110011",
    "1111101101001101",
    "1111101001001011",
    "1111100101011011",
    "1111100001110000",
    "1111011101110011",
    "1111011001010001",
    "1111010100000101",
    "1111001110001111",
    "1111001000000100",
    "1111000010001000",
    "1110111101000100",
    "1110111001011101",
    "1110110111100101",
    "1110110111011111",
    "1110111000110111",
    "1110111011001110",
    "1110111110000111",
    "1111000001001010",
    "1111000100010010",
    "1111000111100010",
    "1111001011010011",
    "1111010000000000",
    "1111010110001011",
    "1111011110001010",
    "1111101000000110",
    "1111110011101101",
    "1111111111100111",
    "1111110010111111",
    "1111100111011111",
    "1111011110001100",
    "1111010111110100",
    "1111010100100101",
    "1111010100011010",
    "1111010110110010",
    "1111011011010100",
    "1111100001100100",
    "1111101001001100",
    "1111110001110110",
    "1111111011000000",
    "1111111100000010",
    "1111110100010000",
    "1111101110100000",
    "1111101011010110",
    "1111101010110110",
    "1111101100011001",
    "1111101110111111",
    "1111110001010110",
    "1111110010010001",
    "1111110000111010",
    "1111101100110111",
    "1111100110001001",
    "1111011101001010",
    "1111010010100110",
    "1111000111010110",
    "1110111100100001",
    "1110110011001011",
    "1110101100010111",
    "1110101000101101",
    "1110101000011010",
    "1110101011000100",
    "1110101111110101",
    "1110110101100010",
    "1110111010111111",
    "1110111111001010",
    "1111000001010101",
    "1111000001001010",
    "1110111110101101",
    "1110111010010100",
    "1110110100100111",
    "1110101110001101",
    "1110100111110101",
    "1110100001111110",
    "1110011101000010",
    "1110011001001100",
    "1110010110011101",
    "1110010100101100",
    "1110010011101100",
    "1110010011011000",
    "1110010011101110",
    "1110010100110011",
    "1110010110101101",
    "1110011001100011",
    "1110011101010111",
    "1110100010000010",
    "1110100111010011",
    "1110101100110111",
    "1110110010010111",
    "1110110111100011",
    "1110111100010110",
    "1111000000110110",
    "1111000101011010",
    "1111001010100000",
    "1111010000110101",
    "1111011000111110",
    "1111100011011000",
    "1111110000000011",
    "1111111110011110",
    "1111110010011001",
    "1111100100000001",
    "1111010111110100",
    "1111001110111010",
    "1111001010000010",
    "1111001001011000",
    "1111001100110000",
    "1111010011111001",
    "1111011110011111",
    "1111101100001010",
    "1111111100001001",
    "1111110010110101",
    "1111100010100100",
    "1111010100110100",
    "1111001010111101",
    "1111000101101001",
    "1111000100011101",
    "1111000110011010",
    "1111001010000100",
    "1111001110010010",
    "1111010010011101",
    "1111010110100010",
    "1111011010101111",
    "1111011111010110",
    "1111100100010111",
    "1111101001011111",
    "1111101110010000",
    "1111110010001001",
    "1111110100111010",
    "1111110110100110",
    "1111110111100100",
    "1111111000011011",
    "1111111001110101",
    "1111111100011110",
    "1111111111000011",
    "1111111000011001",
    "1111101111010111",
    "1111100100001101",
    "1111010111100111",
    "1111001010100010",
    "1110111110000010",
    "1110110011000101",
    "1110101010011000",
    "1110100100010000",
    "1110100000110000",
    "1110011111100100",
    "1110100000011001",
    "1110100010111001",
    "1110100110101111",
    "1110101011101011",
    "1110110001011100",
    "1110110111110101",
    "1110111110101001",
    "1111000101110010",
    "1111001101001111",
    "1111010101001000",
    "1111011101100100",
    "1111100110100000",
    "1111101111100011",
    "1111110111111011",
    "1111111110100010",
    "1111111101101001",
    "1111111101011110",
    "1111111110110011",
    "1111110111101110",
    "1111101110010011",
    "1111100100000011",
    "1111011010101011",
    "1111010011101100",
    "1111010000001101",
    "1111010000101110",
    "1111010100111100",
    "1111011011111111",
    "1111100100011100",
    "1111101100101101",
    "1111110011011111",
    "1111110111110110",
    "1111111001011010",
    "1111111000010010",
    "1111110100111011",
    "1111101111111011",
    "1111101001111010",
    "1111100011011111",
    "1111011101011100",
    "1111011000101100",
    "1111010110010110",
    "1111010111011101",
    "1111011100101011",
    "1111100101110100",
    "1111110001111000",
    "1111111111000110",
    "1111110100100010",
    "1111101010111110",
    "1111100101010101",
    "1111100011111100",
    "1111100110011011",
    "1111101011111000",
    "1111110011010110",
    "1111111100000110",
    "1111111010010101",
    "1111110000010011",
    "1111100101111110",
    "1111011011100110",
    "1111010001100010",
    "1111001000001011",
    "1110111111111000",
    "1110111000111001",
    "1110110011010111",
    "1110101111011001",
    "1110101101000000",
    "1110101100010011",
    "1110101101010110",
    "1110110000001010",
    "1110110100110110",
    "1110111011011011",
    "1111000100001000",
    "1111001111000100",
    "1111011100001110",
    "1111101011010010",
    "1111111011011001",
    "1111110100101011",
    "1111100110010101",
    "1111011010100110",
    "1111010010000011",
    "1111001100011100",
    "1111001001000111",
    "1111000111001011",
    "1111000101111100",
    "1111000101010000",
    "1111000101011010",
    "1111000111000011",
    "1111001010101111",
    "1111010000110110",
    "1111011001010101",
    "1111100011101010",
    "1111101111000101",
    "1111111010100111",
    "1111111010100111",
    "1111110001101001",
    "1111101011001001",
    "1111100111100001",
    "1111100110101100",
    "1111101000000010",
    "1111101010011001",
    "1111101100010011",
    "1111101100001111",
    "1111101001001010",
    "1111100010100001",
    "1111011000011011",
    "1111001011011101",
    "1110111100101101",
    "1110101101100001",
    "1110011111010111",
    "1110010011101100",
    "1110001011101011",
    "1110000111111110",
    "1110001000110100",
    "1110001101110101",
    "1110010110100000",
    "1110100010001000",
    "1110110000001111",
    "1111000000011100",
    "1111010010010100",
    "1111100101001001",
    "1111110111110001",
    "1111110111010010",
    "1111101001101011",
    "1111100000101001",
    "1111011100110000",
    "1111011101110101",
    "1111100011000001",
    "1111101011001101",
    "1111110101010000",
    "1111111111110001",
    "1111110100101111",
    "1111101010011000",
    "1111100001011110",
    "1111011010101111",
    "1111010110101101",
    "1111010101101010",
    "1111010111010011",
    "1111011010111100",
    "1111011111101100",
    "1111100100100111",
    "1111101000110111",
    "1111101011111010",
    "1111101101011110",
    "1111101101100100",
    "1111101100011010",
    "1111101010011001",
    "1111100111111111",
    "1111100101101110",
    "1111100100000001",
    "1111100011001011",
    "1111100011001011",
    "1111100011111001",
    "1111100101001011",
    "1111100110111001",
    "1111101001001101",
    "1111101100100010",
    "1111110001011111",
    "1111111000101111",
    "1111111101010110",
    "1111110001000100",
    "1111100011011100",
    "1111010110000100",
    "1111001010110010",
    "1111000011000110",
    "1110111111111010",
    "1111000001001111",
    "1111000110100111",
    "1111001111010111",
    "1111011011000010",
    "1111101001100010",
    "1111111010111101",
    "1111110000111111",
    "1111011011100101",
    "1111000111000011",
    "1110110110010010",
    "1110101011111010",
    "1110101001011110",
    "1110101110111111",
    "1110111010110111",
    "1111001010101000",
    "1111011011101000",
    "1111101011110000",
    "1111111001110011",
    "1111111010101100",
    "1111110001111100",
    "1111101011111000",
    "1111101000011100",
    "1111100111011011",
    "1111101000011011",
    "1111101010100101",
    "1111101100110111",
    "1111101110001001",
    "1111101101100100",
    "1111101010101111",
    "1111100101111001",
    "1111011111101011",
    "1111011000111010",
    "1111010010010101",
    "1111001100100110",
    "1111000111111111",
    "1111000100101111",
    "1111000010111001",
    "1111000010011010",
    "1111000011001000",
    "1111000100111001",
    "1111000111100000",
    "1111001010110101",
    "1111001110101101",
    "1111010011000101",
    "1111010111110111",
    "1111011100111010",
    "1111100001111001",
    "1111100110011000",
    "1111101001111101",
    "1111101100010011",
    "1111101101010101",
    "1111101101011000",
    "1111101101000111",
    "1111101101011000",
    "1111101110111110",
    "1111110010010101",
    "1111110111010110",
    "1111111101011001",
    "1111111100011010",
    "1111110111001010",
    "1111110011100101",
    "1111110010000110",
    "1111110010101110",
    "1111110101001000",
    "1111111000111000",
    "1111111101101000",
    "1111111100111010",
    "1111110111000011",
    "1111110001001001",
    "1111101011101010",
    "1111100111010010",
    "1111100100110001",
    "1111100100110001",
    "1111100111101011",
    "1111101101011101",
    "1111110101101110",
    "1111111111101010",
    "1111110101100101",
    "1111101011001001",
    "1111100001111000",
    "1111011010100110",
    "1111010101111011",
    "1111010100001000",
    "1111010101010011",
    "1111011001001110",
    "1111011111010010",
    "1111100110110000",
    "1111101110100101",
    "1111110101101111",
    "1111111011010111",
    "1111111110111000",
    "1111111111110110",
    "1111111111011110",
    "1111111101101101",
    "1111111011101111",
    "1111111010011101",
    "1111111010100001",
    "1111111100010000",
    "1111111111110100",
    "1111111010101110",
    "1111110011011001",
    "1111101010000100",
    "1111011110111011",
    "1111010010100110",
    "1111000110001001",
    "1110111010111111",
    "1110110010011101",
    "1110101101100110",
    "1110101100110010",
    "1110101111111000",
    "1110110110011011",
    "1110111111111010",
    "1111001011110111",
    "1111011001111010",
    "1111101001100010",
    "1111111001110101",
    "1111110110010100",
    "1111101000010001",
    "1111011101000000",
    "1111010101000101",
    "1111010000010111",
    "1111001110010111",
    "1111001110010100",
    "1111001111100100",
    "1111010001110100",
    "1111010101000011",
    "1111011001011110",
    "1111011111010111",
    "1111100110111011",
    "1111110000010101",
    "1111111011101110",
    "1111110110111101",
    "1111101000001100",
    "1111011000111010",
    "1111001010110010",
    "1110111111101110",
    "1110111001100010",
    "1110111001010011",
    "1110111111000111",
    "1111001001110101",
    "1111010111011010",
    "1111100101011010",
    "1111110001100111",
    "1111111010011011",
    "1111111111001100",
    "1111111111111001",
    "1111111101111001",
    "1111111001110111",
    "1111110101010001",
    "1111110001010101",
    "1111101111000001",
    "1111101111000010",
    "1111110001101101",
    "1111110110111110",
    "1111111110001111",
    "1111111001010111",
    "1111110001000111",
    "1111101010000101",
    "1111100101001001",
    "1111100010111000",
    "1111100011011100",
    "1111100110101001",
    "1111101100001100",
    "1111110011100110",
    "1111111100011010",
    "1111111001110000",
    "1111101111011110",
    "1111100101001101",
    "1111011011100011",
    "1111010011000000",
    "1111001011111010",
    "1111000110010101",
    "1111000010000110",
    "1110111110111010",
    "1110111100011001",
    "1110111010010110",
    "1110111000110000",
    "1110110111101111",
    "1110110111010110",
    "1110110111101111",
    "1110111000110100",
    "1110111010011000",
    "1110111100010100",
    "1110111110100011",
    "1111000001001101",
    "1111000100101010",
    "1111001001100010",
    "1111010000011010",
    "1111011001110101",
    "1111100101111100",
    "1111110100010101",
    "1111111100000011",
    "1111101100101111",
    "1111011111011001",
    "1111010101011011",
    "1111001111110000",
    "1111001110011111",
    "1111010001000101",
    "1111010110100010",
    "1111011101110011",
    "1111100101111110",
    "1111101110011101",
    "1111110111000000",
    "1111111111011101",
    "1111111000010001",
    "1111110000011111",
    "1111101001100110",
    "1111100100000000",
    "1111100000000010",
    "1111011101110111",
    "1111011101010100",
    "1111011110000000",
    "1111011111011010",
    "1111100000111110",
    "1111100010010010",
    "1111100011000001",
    "1111100011001011",
    "1111100010111101",
    "1111100010101011",
    "1111100010110011",
    "1111100011110011",
    "1111100110000011",
    "1111101001111000",
    "1111101111100111",
    "1111110111011000",
    "1111111110110100",
    "1111110011100001",
    "1111100111100011",
    "1111011100000100",
    "1111010010010101",
    "1111001011010110",
    "1111000111110001",
    "1111000111101100",
    "1111001010110101",
    "1111010000101011",
    "1111011000101000",
    "1111100010010100",
    "1111101101010101",
    "1111111001011011",
    "1111111001110011",
    "1111101100111110",
    "1111100000110000",
    "1111010101110100",
    "1111001100101011",
    "1111000101100101",
    "1111000000011111",
    "1110111101000000",
    "1110111010110100",
    "1110111001100000",
    "1110111000110111",
    "1110111000101101",
    "1110111001000100",
    "1110111001111101",
    "1110111011011101",
    "1110111101100001",
    "1111000000000111",
    "1111000010111101",
    "1111000101110010",
    "1111001000011000",
    "1111001010100011",
    "1111001100011001",
    "1111001110000010",
    "1111001111110001",
    "1111010001111000",
    "1111010100011101",
    "1111010111011111",
    "1111011010111000",
    "1111011110011110",
    "1111100010000110",
    "1111100101110010",
    "1111101001101101",
    "1111101110001011",
    "1111110011100001",
    "1111111001111011",
    "1111111110101101",
    "1111110110110101",
    "1111101111000111",
    "1111101000010010",
    "1111100010111011",
    "1111011111011001",
    "1111011101101011",
    "1111011101011100",
    "1111011101111111",
    "1111011110011110",
    "1111011110000000",
    "1111011011110000",
    "1111010111001110",
    "1111010000010010",
    "1111000111010101",
    "1110111101001001",
    "1110110010101111",
    "1110101001010011",
    "1110100001110001",
    "1110011100111010",
    "1110011010111100",
    "1110011011101111",
    "1110011110111000",
    "1110100011101100",
    "1110101001011101",
    "1110101111100001",
    "1110110101010011",
    "1110111010011011",
    "1110111110101110",
    "1111000010010010",
    "1111000101011000",
    "1111001000011110",
    "1111001100000001",
    "1111010000011010",
    "1111010101111001",
    "1111011100010111",
    "1111100011100111",
    "1111101011001110",
    "1111110010110000",
    "1111111001110101",
    "1111111111110011",
    "1111111010011001",
    "1111110110000100",
    "1111110010111100",
    "1111110001000110",
    "1111110000110001",
    "1111110010001000",
    "1111110101011000",
    "1111111010101011",
    "1111111101110011",
    "1111110100000100",
    "1111101000001101",
    "1111011010100011",
    "1111001011110010",
    "1110111100111100",
    "1110101111010111",
    "1110100100010111",
    "1110011100111111",
    "1110011001101111",
    "1110011010011001",
    "1110011110001100",
    "1110100011111000",
    "1110101010000100",
    "1110101111011110",
    "1110110011001011",
    "1110110100100100",
    "1110110011100010",
    "1110110000010100",
    "1110101011010110",
    "1110100101011101",
    "1110011111011110",
    "1110011010010001",
    "1110010110101010",
    "1110010101001000",
    "1110010110000001",
    "1110011001010101",
    "1110011110111111",
    "1110100110110100",
    "1110110000101110",
    "1110111100100110",
    "1111001010010011",
    "1111011001010001",
    "1111101000101101",
    "1111110111010110",
    "1111111100000101",
    "1111110010101110",
    "1111101101000111",
    "1111101011001000",
    "1111101100000011",
    "1111101110110101",
    "1111110010011010",
    "1111110101111110",
    "1111111001000010",
    "1111111011011100",
    "1111111101001100",
    "1111111110010010",
    "1111111110101011",
    "1111111110010010",
    "1111111101000100",
    "1111111011000001",
    "1111111000010010",
    "1111110101000001",
    "1111110001011011",
    "1111101101100100",
    "1111101001100110",
    "1111100101100000",
    "1111100001011001",
    "1111011101010111",
    "1111011001101011",
    "1111010110101100",
    "1111010100110111",
    "1111010100110100",
    "1111010111001001",
    "1111011100100101",
    "1111100101100000",
    "1111110010000101",
    "1111111110010000",
    "1111101100111000",
    "1111011011100101",
    "1111001100010011",
    "1111000000101110",
    "1110111001110000",
    "1110110111100101",
    "1110111001100101",
    "1110111110110101",
    "1111000110010011",
    "1111001111000111",
    "1111011000010001",
    "1111100000101100",
    "1111100111000010",
    "1111101001110110",
    "1111101000001011",
    "1111100001110011",
    "1111010111101010",
    "1111001011101000",
    "1111000000001101",
    "1110110111101100",
    "1110110011101001",
    "1110110100100100",
    "1110111001110101",
    "1111000010010100",
    "1111001100101000",
    "1111010111101101",
    "1111100010111000",
    "1111101101101110",
    "1111111000000011",
    "1111111110010111",
    "1111110101111110",
    "1111101111001010",
    "1111101010010010",
    "1111100111100100",
    "1111100110111001",
    "1111100111111111",
    "1111101010011010",
    "1111101101101100",
    "1111110001011001",
    "1111110101001010",
    "1111111000101011",
    "1111111011101010",
    "1111111101111000",
    "1111111111001000",
    "1111111111010010",
    "1111111110010011",
    "1111111100001110",
    "1111111001000110",
    "1111110101000100",
    "1111110000010000",
    "1111101010110111",
    "1111100101001101",
    "1111011111100110",
    "1111011010011001",
    "1111010101111100",
    "1111010010010111",
    "1111001111101110",
    "1111001101111011",
    "1111001100111010",
    "1111001100101000",
    "1111001101000111",
    "1111001110100011",
    "1111010001000000",
    "1111010100100100",
    "1111011001000110",
    "1111011110001100",
    "1111100011010101",
    "1111100111111111",
    "1111101011101000",
    "1111101101111011",
    "1111101110101110",
    "1111101110000011",
    "1111101100000111",
    "1111101001001010",
    "1111100101011011",
    "1111100001010010",
    "1111011101000010",
    "1111011001000100",
    "1111010101110111",
    "1111010011111100",
    "1111010011110110",
    "1111010101111001",
    "1111011010001100",
    "1111100000011100",
    "1111101000000010",
    "1111110000000111",
    "1111110111101010",
    "1111111101110100",
    "1111111101111110",
    "1111111100000011",
    "1111111100010011",
    "1111111110011011",
    "1111111101111100",
    "1111111001010000",
    "1111110011101100",
    "1111101101010011",
    "1111100110000011",
    "1111011101110111",
    "1111010100110001",
    "1111001011000001",
    "1111000001000000",
    "1110110111010110",
    "1110101110101110",
    "1110100111101100",
    "1110100010100001",
    "1110011111010001",
    "1110011101101000",
    "1110011101000111",
    "1110011101000111",
    "1110011101000100",
    "1110011100101000",
    "1110011011101010",
    "1110011010001001",
    "1110011000010101",
    "1110010110100000",
    "1110010101000000",
    "1110010100000101",
    "1110010011111110",
    "1110010100110011",
    "1110010110100111",
    "1110011001010110",
    "1110011100110011",
    "1110100000110000",
    "1110100100110100",
    "1110101000101111",
    "1110101100010111",
    "1110101111101011",
    "1110110010111001",
    "1110110110010110",
    "1110111010100101",
    "1110111111111000",
    "1111000110011111",
    "1111001110001101",
    "1111010110100101",
    "1111011110110000",
    "1111100101101111",
    "1111101010011001",
    "1111101011110011",
    "1111101001010101",
    "1111100010111001",
    "1111011001010001",
    "1111001101111010",
    "1111000010110100",
    "1110111010001001",
    "1110110101011111",
    "1110110101110001",
    "1110111011000001",
    "1111000100100111",
    "1111010001101011",
    "1111100001010111",
    "1111110010111100",
    "1111111010011010",
    "1111101000000100",
    "1111010111101101",
    "1111001011010001",
    "1111000100011101",
    "1111000100001110",
    "1111001010100101",
    "1111010110100010",
    "1111100110010011",
    "1111110111101101",
    "1111110111010010",
    "1111101000100011",
    "1111011101001110",
    "1111010101111001",
    "1111010010100010",
    "1111010010101110",
    "1111010101100111",
    "1111011010011000",
    "1111100000010100",
    "1111100110111010",
    "1111101101110111",
    "1111110101000100",
    "1111111100011000",
    "1111111100010110",
    "1111110101100100",
    "1111101111110010",
    "1111101011100010",
    "1111101001001100",
    "1111101000110110",
    "1111101010001100",
    "1111101100101100",
    "1111101111101010",
    "1111110010011000",
    "1111110100001111",
    "1111110100110100",
    "1111110011111010",
    "1111110001100110",
    "1111101110001011",
    "1111101010000111",
    "1111100101111110",
    "1111100010010000",
    "1111011111011001",
    "1111011101100000",
    "1111011100011100",
    "1111011011110111",
    "1111011011001001",
    "1111011001101011",
    "1111010110111111",
    "1111010010110110",
    "1111001101011100",
    "1111000111010110",
    "1111000001100001",
    "1110111100110101",
    "1110111010001100",
    "1110111010001100",
    "1110111101000000",
    "1111000010011111",
    "1111001010001111",
    "1111010011110001",
    "1111011110011100",
    "1111101001100001",
    "1111110100000010",
    "1111111100110110",
    "1111111101000100",
    "1111111010100001",
    "1111111011101100",
    "1111111111111000",
    "1111111001001011",
    "1111110001010011",
    "1111101001001110",
    "1111100001100001",
    "1111011010010001",
    "1111010011010111",
    "1111001100101010",
    "1111000110001011",
    "1111000000010100",
    "1110111011101101",
    "1110111000111010",
    "1110111000010110",
    "1110111010000010",
    "1110111101101000",
    "1111000010011100",
    "1111000111101010",
    "1111001100100001",
    "1111010000100011",
    "1111010011100010",
    "1111010101101010",
    "1111010111010011",
    "1111011000111010",
    "1111011011000010",
    "1111011101111101",
    "1111100001111011",
    "1111100111000101",
    "1111101101011101",
    "1111110100111101",
    "1111111101010010",
    "1111111010000011",
    "1111110001110100",
    "1111101010110000",
    "1111100101100010",
    "1111100010100010",
    "1111100001111101",
    "1111100011101010",
    "1111100111011010",
    "1111101100110110",
    "1111110011101000",
    "1111111011011101",
    "1111111011111011",
    "1111110010111000",
    "1111101001100110",
    "1111100000010001",
    "1111010111001000",
    "1111001110010010",
    "1111000110000011",
    "1110111110101000",
    "1110111000011110",
    "1110110100000110",
    "1110110010000110",
    "1110110011000110",
    "1110110111110010",
    "1111000000101100",
    "1111001110000100",
    "1111011111010111",
    "1111110011000100",
    "1111111001001101",
    "1111101000010001",
    "1111011100011110",
    "1111010111000110",
    "1111011000001000",
    "1111011110010010",
    "1111100111110010",
    "1111110010111010",
    "1111111110110000",
    "1111110100111011",
    "1111101000001011",
    "1111011011001111",
    "1111001111001000",
    "1111000101011000",
    "1110111111100100",
    "1110111110110101",
    "1111000011001000",
    "1111001011010001",
    "1111010101001101",
    "1111011110100110",
    "1111100101011111",
    "1111101000101010",
    "1111100111110000",
    "1111100011000000",
    "1111011011000111",
    "1111010001001100",
    "1111000110011010",
    "1110111100000100",
    "1110110011011100",
    "1110101101100100",
    "1110101011010011",
    "1110101101000111",
    "1110110011010000",
    "1110111101110011",
    "1111001100100001",
    "1111011110111000",
    "1111110011110101",
    "1111110110000111",
    "1111100000111101",
    "1111001110011100",
    "1110111111111111",
    "1110110110000001",
    "1110110000001100",
    "1110101101011100",
    "1110101100100110",
    "1110101100101011",
    "1110101101010001",
    "1110101110011011",
    "1110110000011100",
    "1110110011011111",
    "1110110111011101",
    "1110111100000001",
    "1111000000101011",
    "1111000101000101",
    "1111001001001001",
    "1111001101001100",
    "1111010001101110",
    "1111010111011000",
    "1111011110101001",
    "1111100111111101",
    "1111110011100101",
    "1111111110010100",
    "1111101110000010",
    "1111011100011110",
    "1111001011000111",
    "1110111011110101",
    "1110110000010010",
    "1110101001100011",
    "1110100111101100",
    "1110101001110111",
    "1110101110101000",
    "1110110100100010",
    "1110111010100011",
    "1111000000010010",
    "1111000101110110",
    "1111001011100011",
    "1111010001101001",
    "1111011000000011",
    "1111011110011110",
    "1111100100100010",
    "1111101001111100",
    "1111101110101001",
    "1111110010111110",
    "1111110111010100",
    "1111111100000001",
    "1111111110110011",
    "1111111001011111",
    "1111110100011110",
    "1111110000001111",
    "1111101101001010",
    "1111101011011011",
    "1111101010111010",
    "1111101011010011",
    "1111101100001100",
    "1111101101001111",
    "1111101110001110",
    "1111101111000101",
    "1111101111110100",
    "1111110000100001",
    "1111110001001101",
    "1111110001110101",
    "1111110010001110",
    "1111110010000101",
    "1111110001000110",
    "1111101111000001",
    "1111101011101001",
    "1111100111000011",
    "1111100001011010",
    "1111011011001110",
    "1111010100111100",
    "1111001111000111",
    "1111001010001001",
    "1111000110010101",
    "1111000011110110",
    "1111000010101110",
    "1111000011000000",
    "1111000100101100",
    "1111000111110111",
    "1111001100100101",
    "1111010011000011",
    "1111011011011011",
    "1111100101110111",
    "1111110010011101",
    "1111111111000100",
    "1111101111011001",
    "1111011111011110",
    "1111010000100001",
    "1111000011101100",
    "1110111001110100",
    "1110110011010101",
    "1110110000000111",
    "1110101111110000",
    "1110110001101100",
    "1110110101011000",
    "1110111010011001",
    "1111000000011100",
    "1111000111001000",
    "1111001101111010",
    "1111010100000001",
    "1111011000101000",
    "1111011011000100",
    "1111011011000010",
    "1111011000111111",
    "1111010101111110",
    "1111010011100001",
    "1111010011010000",
    "1111010110011111",
    "1111011101111010",
    "1111101001100011",
    "1111111000101001",
    "1111110110000011",
    "1111100100010010",
    "1111010011110001",
    "1111000110001000",
    "1110111100100001",
    "1110110111100111",
    "1110110111010001",
    "1110111010111010",
    "1111000001011010",
    "1111001001100010",
    "1111010010000011",
    "1111011010000010",
    "1111100000111000",
    "1111100110001110",
    "1111101010000110",
    "1111101100101010",
    "1111101110001110",
    "1111101111010000",
    "1111110000010010",
    "1111110001110010",
    "1111110100010001",
    "1111111000000001",
    "1111111101000111",
    "1111111100101010",
    "1111110101111011",
    "1111101111011000",
    "1111101001111000",
    "1111100110000100",
    "1111100100011101",
    "1111100101001000",
    "1111100111111001",
    "1111101100100001",
    "1111110010101100",
    "1111111010010000",
    "1111111100110010",
    "1111110010100011",
    "1111100111010101",
    "1111011011110011",
    "1111010001001100",
    "1111001000110111",
    "1111000100010000",
    "1111000100010111",
    "1111001001101000",
    "1111010011111000",
    "1111100010000110",
    "1111110010101110",
    "1111111100000110",
    "1111101100011001",
    "1111011111101011",
    "1111010110111011",
    "1111010010010111",
    "1111010001100110",
    "1111010011101100",
    "1111010111100010",
    "1111011100000100",
    "1111100000011110",
    "1111100100001011",
    "1111100110110101",
    "1111101000010001",
    "1111101000011100",
    "1111100111011100",
    "1111100101100000",
    "1111100011000101",
    "1111100000101110",
    "1111011111000100",
    "1111011110101000",
    "1111011111110011",
    "1111100010101111",
    "1111100111011110",
    "1111101101111011",
    "1111110110001011",
    "1111111111101010",
    "1111110011100110",
    "1111100101110001",
    "1111010110110110",
    "1111001000000100",
    "1110111011000100",
    "1110110001100110",
    "1110101101000100",
    "1110101110001010",
    "1110110100110100",
    "1111000000001000",
    "1111001110101101",
    "1111011110110001",
    "1111101110110001",
    "1111111101010101",
    "1111110110011101",
    "1111101101001110",
    "1111100111000110",
    "1111100011111100",
    "1111100011011100",
    "1111100101000011",
    "1111101000010110",
    "1111101100111010",
    "1111110010010011",
    "1111111000010001",
    "1111111110100011",
    "1111111010111110",
    "1111110100011110",
    "1111101101111111",
    "1111100111100000",
    "1111100001000011",
    "1111011010100110",
    "1111010100010111",
    "1111001110100110",
    "1111001001110101",
    "1111000110011111",
    "1111000100110111",
    "1111000100111011",
    "1111000110010010",
    "1111001000000100",
    "1111001001010001",
    "1111001000110100",
    "1111000101110100",
    "1110111111110110",
    "1110110111001110",
    "1110101100110010",
    "1110100010000000",
    "1110011000101101",
    "1110010010011111",
    "1110010000100100",
    "1110010011011100",
    "1110011010111000",
    "1110100110001001",
    "1110110100001011",
    "1111000011110100",
    "1111010100000110",
    "1111100100000110",
    "1111110010111100",
    "1111111111101010",
    "1111110110101010",
    "1111110000111100",
    "1111101111101010",
    "1111110010110000",
    "1111111001101100",
    "1111111100100110",
    "1111110001100101",
    "1111100110101001",
    "1111011101000010",
    "1111010101101001",
    "1111010000111101",
    "1111001111000000",
    "1111001111100011",
    "1111010001111000",
    "1111010101010011",
    "1111011000111111",
    "1111011100001111",
    "1111011110100110",
    "1111011111111010",
    "1111100000001100",
    "1111011111101100",
    "1111011110110101",
    "1111011101111000",
    "1111011101001001",
    "1111011100110010",
    "1111011100111000",
    "1111011101100001",
    "1111011110101110",
    "1111100000011100",
    "1111100010101001",
    "1111100101001110",
    "1111100111111110",
    "1111101010101010",
    "1111101101000001",
    "1111101110110101",
    "1111101111111101",
    "1111110000010010",
    "1111101111111011",
    "1111101111000001",
    "1111101101111000",
    "1111101100110110",
    "1111101100010001",
    "1111101100011110",
    "1111101101110000",
    "1111110000010100",
    "1111110100001101",
    "1111111001001101",
    "1111111110110100",
    "1111111011110110",
    "1111111000000101",
    "1111110111000110",
    "1111111001111110",
    "1111111110110110",
    "1111110011111101",
    "1111100110110010",
    "1111011001011001",
    "1111001101111101",
    "1111000110001000",
    "1111000010110100",
    "1111000011111100",
    "1111001000101101",
    "1111001111110011",
    "1111010111110010",
    "1111011111100100",
    "1111100110010101",
    "1111101011111001",
    "1111110000110010",
    "1111110110000110",
    "1111111101000100",
    "1111111001011111",
    "1111101101110000",
    "1111100000110000",
    "1111010100010011",
    "1111001010011110",
    "1111000100111100",
    "1111000100011100",
    "1111001000011101",
    "1111001111101001",
    "1111011000000100",
    "1111011111111101",
    "1111100101110111",
    "1111101001001010",
    "1111101001101101",
    "1111101000000000",
    "1111100100101110",
    "1111100000101011",
    "1111011100101011",
    "1111011001100000",
    "1111010111110111",
    "1111011000010110",
    "1111011011001110",
    "1111100000001101",
    "1111100110110001",
    "1111101101110111",
    "1111110100011111",
    "1111111001101010",
    "1111111100110101",
    "1111111101110101",
    "1111111100111101",
    "1111111010110000",
    "1111110111110101",
    "1111110100101010",
    "1111110001100010",
    "1111101110100100",
    "1111101011100111",
    "1111101000100010",
    "1111100100111100",
    "1111100000100011",
    "1111011010111000",
    "1111010011101110",
    "1111001010111111",
    "1111000000111001",
    "1110110110000011",
    "1110101011011011",
    "1110100010001111",
    "1110011011101101",
    "1110011000111110",
    "1110011010101101",
    "1110100001000011",
    "1110101011011110",
    "1110111000101111",
    "1111000111000011",
    "1111010100010011",
    "1111011110011111",
    "1111100100010000",
    "1111100100110111",
    "1111100000101001",
    "1111011000010110",
    "1111001101000100",
    "1110111111110000",
    "1110110001010100",
    "1110100010101001",
    "1110010100110011",
    "1110001000111100",
    "1110000000000111",
    "1101111011000010",
    "1101111001111100",
    "1101111100011001",
    "1110000001100110",
    "1110001000100011",
    "1110010000010111",
    "1110011000010011",
    "1110011111110110",
    "1110100110100101",
    "1110101100001100",
    "1110110000010001",
    "1110110010100001",
    "1110110010110011",
    "1110110001010100",
    "1110101110100011",
    "1110101011010100",
    "1110101000011101",
    "1110100110101100",
    "1110100110101100",
    "1110101000110111",
    "1110101101011001",
    "1110110100011100",
    "1110111101111010",
    "1111001001101111",
    "1111010111110001",
    "1111100111101100",
    "1111111000111110",
    "1111110101010001",
    "1111100100011000",
    "1111010101101111",
    "1111001010100011",
    "1111000011011111",
    "1111000000100110",
    "1111000001001101",
    "1111000100001010",
    "1111001000001110",
    "1111001100011100",
    "1111010000011001",
    "1111010100000110",
    "1111011000000100",
    "1111011101000101",
    "1111100011111011",
    "1111101101001000",
    "1111111001000000",
    "1111111000101001",
    "1111101000100101",
    "1111011000000110",
    "1111001001000110",
    "1110111101100011",
    "1110110111000110",
    "1110110110011011",
    "1110111011001010",
    "1111000011111011",
    "1111001110101011",
    "1111011001100000",
    "1111100010111110",
    "1111101010011001",
    "1111101111101010",
    "1111110011000010",
    "1111110100110111",
    "1111110101010111",
    "1111110100100100",
    "1111110010100101",
    "1111101111100101",
    "1111101100000000",
    "1111101000011011",
    "1111100101100000",
    "1111100011110110",
    "1111100011101111",
    "1111100101010111",
    "1111101000110001",
    "1111101110000001",
    "1111110101000100",
    "1111111101100111",
    "1111111000111110",
    "1111101111110000",
    "1111100111111011",
    "1111100010100110",
    "1111100000100100",
    "1111100010000101",
    "1111100110110001",
    "1111101101101011",
    "1111110101100011",
    "1111111101000101",
    "1111111100111001",
    "1111111001010000",
    "1111111000100100",
    "1111111011000000",
    "1111111111011000",
    "1111110110111000",
    "1111101011111010",
    "1111011111010001",
    "1111010010000000",
    "1111000101011000",
    "1110111010101011",
    "1110110010111001",
    "1110101110101101",
    "1110101110010001",
    "1110110001010100",
    "1110110111010101",
    "1110111111011111",
    "1111001000111100",
    "1111010010111001",
    "1111011100100110",
    "1111100101100111",
    "1111101101101100",
    "1111110100110110",
    "1111111011010101",
    "1111111110100011",
    "1111111000101011",
    "1111110010111110",
    "1111101101101100",
    "1111101001001011",
    "1111100101110110",
    "1111100011111110",
    "1111100011110001",
    "1111100101010000",
    "1111101000011011",
    "1111101101010011",
    "1111110011111001",
    "1111111100001011",
    "1111111010001001",
    "1111101111110110",
    "1111100110000110",
    "1111011110010111",
    "1111011001111111",
    "1111011001111100",
    "1111011110001100",
    "1111100101110010",
    "1111101110111001",
    "1111110111010010",
    "1111111100111100",
    "1111111110011111",
    "1111111011100001",
    "1111110100100001",
    "1111101010100110",
    "1111011111000100",
    "1111010011001000",
    "1111000111110111",
    "1110111110000100",
    "1110110110011010",
    "1110110001100110",
    "1110110000000011",
    "1110110010000011",
    "1110110111011010",
    "1110111111100011",
    "1111001001100111",
    "1111010100100000",
    "1111011111010010",
    "1111101001001001",
    "1111110001100001",
    "1111111000001110",
    "1111111101010001",
    "1111111111000101",
    "1111111100101011",
    "1111111011010100",
    "1111111010110111",
    "1111111011010001",
    "1111111100100001",
    "1111111110100110",
    "1111111110011111",
    "1111111010111100",
    "1111110110110111",
    "1111110010011011",
    "1111101101110100",
    "1111101001000100",
    "1111100100001010",
    "1111011110111010",
    "1111011000111110",
    "1111010001111011",
    "1111001001011110",
    "1110111111101000",
    "1110110100111001",
    "1110101010010100",
    "1110100001001101",
    "1110011010110010",
    "1110010111110010",
    "1110011000010011",
    "1110011011101011",
    "1110100000111011",
    "1110100110110111",
    "1110101100100101",
    "1110110001011100",
    "1110110101001001",
    "1110110111100111",
    "1110111000101100",
    "1110111000010110",
    "1110110110101010",
    "1110110011110001",
    "1110110000000111",
    "1110101100010100",
    "1110101001000100",
    "1110100110111100",
    "1110100110010110",
    "1110100111010101",
    "1110101001101101",
    "1110101101001111",
    "1110110001101001",
    "1110110110110010",
    "1110111100100001",
    "1111000010110001",
    "1111001001011000",
    "1111010000001000",
    "1111010110110110",
    "1111011101001010",
    "1111100010111001",
    "1111100111111100",
    "1111101100010000",
    "1111110000000011",
    "1111110011100110",
    "1111110111010101",
    "1111111011100100",
    "1111111111011000",
    "1111111001100100",
    "1111110011001011",
    "1111101100101100",
    "1111100110101101",
    "1111100001110001",
    "1111011110011100",
    "1111011101000000",
    "1111011101100100",
    "1111100000000111",
    "1111100100010101",
    "1111101001111011",
    "1111110000011001",
    "1111110111001101",
    "1111111101110000",
    "1111111100010110",
    "1111110111011101",
    "1111110011100111",
    "1111110000101010",
    "1111101110010001",
    "1111101100000100",
    "1111101001110000",
    "1111100111000111",
    "1111100100001110",
    "1111100001010101",
    "1111011110111010",
    "1111011101011110",
    "1111011101101000",
    "1111011111111011",
    "1111100100110001",
    "1111101100011000",
    "1111110110101001",
    "1111111100111001",
    "1111101111001110",
    "1111100001011110",
    "1111010100111011",
    "1111001010101000",
    "1111000011011000",
    "1110111111100100",
    "1110111111001101",
    "1111000010001011",
    "1111001000001110",
    "1111010000110011",
    "1111011010111010",
    "1111100101000000",
    "1111101101000110",
    "1111110001010100",
    "1111110000001101",
    "1111101001001100",
    "1111011100101110",
    "1111001100010001",
    "1110111010000001",
    "1110101000011011",
    "1110011001110101",
    "1110001111110110",
    "1110001011001111",
    "1110001011111101",
    "1110010001001010",
    "1110011001100010",
    "1110100011101010",
    "1110101110011011",
    "1110111000111001",
    "1111000010100010",
    "1111001011000111",
    "1111010010100010",
    "1111011000111001",
    "1111011110010001",
    "1111100010101110",
    "1111100110011011",
    "1111101001011000",
    "1111101011110000",
    "1111101101100111",
    "1111101111000110",
    "1111110000001110",
    "1111110001000001",
    "1111110001100010",
    "1111110001111011",
    "1111110010011010",
    "1111110011010110",
    "1111110101000101",
    "1111110111111011",
    "1111111100000110",
    "1111111110011000",
    "1111110111110101",
    "1111110000101010",
    "1111101001011000",
    "1111100010011100",
    "1111011100000101",
    "1111010110011010",
    "1111010001010010",
    "1111001100100011",
    "1111001000000100",
    "1111000011111001",
    "1111000000001100",
    "1110111101001010",
    "1110111011000111",
    "1110111010011000",
    "1110111011000100",
    "1110111101010111",
    "1111000001001111",
    "1111000110100101",
    "1111001101001100",
    "1111010100110100",
    "1111011101000100",
    "1111100101100010",
    "1111101101110011",
    "1111110101011001",
    "1111111011111111",
    "1111111110100110",
    "1111111010011110",
    "1111110111011101",
    "1111110101001011",
    "1111110011001001",
    "1111110000110011",
    "1111101101101101",
    "1111101001100001",
    "1111100100000110",
    "1111011101011110",
    "1111010101101111",
    "1111001101010010",
    "1111000100101010",
    "1110111100100101",
    "1110110101110010",
    "1110110001000000",
    "1110101110101000",
    "1110101110101110",
    "1110110001001101",
    "1110110101101111",
    "1110111100000100",
    "1111000100000101",
    "1111001101100110",
    "1111011000010110",
    "1111100011110011",
    "1111101111000110",
    "1111111001010101",
    "1111111110010111",
    "1111111000101011",
    "1111110101101110",
    "1111110101010001",
    "1111110110110001",
    "1111111001100101",
    "1111111101001011",
    "1111111110110000",
    "1111111010100010",
    "1111110110010000",
    "1111110010000011",
    "1111101110000111",
    "1111101010101100",
    "1111101000001000",
    "1111100110101011",
    "1111100110100100",
    "1111100111110111",
    "1111101010100001",
    "1111101110010010",
    "1111110010111010",
    "1111111000001000",
    "1111111101101001",
    "1111111100110001",
    "1111110111011100",
    "1111110010101100",
    "1111101110110111",
    "1111101100010011",
    "1111101011010001",
    "1111101011111100",
    "1111101110011011",
    "1111110010110101",
    "1111111001010000",
    "1111111110001000",
    "1111110011100110",
    "1111100111110101",
    "1111011100000111",
    "1111010010001000",
    "1111001011100110",
    "1111001001101010",
    "1111001100101110",
    "1111010100001011",
    "1111011110011100",
    "1111101001100001",
    "1111110011001011",
    "1111111001100001",
    "1111111011001011",
    "1111110111011110",
    "1111101110011000",
    "1111100000101001",
    "1111001111101000",
    "1110111101010010",
    "1110101011110010",
    "1110011101000111",
    "1110010010101111",
    "1110001101011001",
    "1110001100111000",
    "1110010000010101",
    "1110010110101100",
    "1110011110110101",
    "1110100111111111",
    "1110110001101011",
    "1110111011011110",
    "1111000101000110",
    "1111001110010010",
    "1111010110110111",
    "1111011110110011",
    "1111100110010110",
    "1111101101111111",
    "1111110110001101",
    "1111111111010101",
    "1111110110110000",
    "1111101100110000",
    "1111100011101001",
    "1111011100010110",
    "1111010111100000",
    "1111010101000011",
    "1111010100011111",
    "1111010100111001",
    "1111010101011000",
    "1111010101010011",
    "1111010100011000",
    "1111010010101111",
    "1111010000110001",
    "1111001110111101",
    "1111001101101101",
    "1111001101011001",
    "1111001110000111",
    "1111001111110001",
    "1111010010000110",
    "1111010100110001",
    "1111010111011000",
    "1111011001101000",
    "1111011011011000",
    "1111011100110010",
    "1111011110001101",
    "1111100000010010",
    "1111100011101110",
    "1111101001000110",
    "1111110000111000",
    "1111111011000010",
    "1111111000111111",
    "1111101100100000",
    "1111100001000011",
    "1111011000010001",
    "1111010011011010",
    "1111010010111110",
    "1111010110101100",
    "1111011101100001",
    "1111100110010010",
    "1111101111100111",
    "1111111000100000",
    "1111111111110100",
    "1111111010000110",
    "1111110110111010",
    "1111110110111001",
    "1111111010100111",
    "1111111101101000",
    "1111110010001010",
    "1111100011111110",
    "1111010100101010",
    "1111000110001000",
    "1110111010000001",
    "1110110001011110",
    "1110101100101101",
    "1110101011010001",
    "1110101100011110",
    "1110101111100100",
    "1110110100010011",
    "1110111010110000",
    "1111000011010011",
    "1111001110010110",
    "1111011011111010",
    "1111101011011100",
    "1111111011110110",
    "1111110100011010",
    "1111100110111110",
    "1111011101000111",
    "1111010111100010",
    "1111010110010010",
    "1111011000101111",
    "1111011101111000",
    "1111100100010101",
    "1111101010101010",
    "1111101111100100",
    "1111110010010001",
    "1111110010100001",
    "1111110000101010",
    "1111101101011011",
    "1111101001100110",
    "1111100101101111",
    "1111100010000101",
    "1111011110101011",
    "1111011011100001",
    "1111011000110101",
    "1111010111000001",
    "1111010110100111",
    "1111011000001001",
    "1111011011111101",
    "1111100010001010",
    "1111101010100001",
    "1111110100101001",
    "1111111111111101",
    "1111110100000111",
    "1111101000010110",
    "1111011101011100",
    "1111010100001010",
    "1111001101001110",
    "1111001001010000",
    "1111001000101101",
    "1111001011110111",
    "1111010010101110",
    "1111011101010010",
    "1111101011100111",
    "1111111101101000",
    "1111101101001001",
    "1111010110001000",
    "1110111111011110",
    "1110101100000001",
    "1110011110011011",
    "1110011000100010",
    "1110011010111100",
    "1110100100110111",
    "1110110100011010",
    "1111000111001000",
    "1111011010011110",
    "1111101100001101",
    "1111111010100000",
    "1111111011110101",
    "1111110111011101",
    "1111111000001100",
    "1111111101001111",
    "1111111010101110",
    "1111110001011010",
    "1111101000011100",
    "1111100001010000",
    "1111011100110000",
    "1111011011010110",
    "1111011100111100",
    "1111100001000011",
    "1111100111001100",
    "1111101110101101",
    "1111110110111101",
    "1111111111010000",
    "1111111001001011",
    "1111110011000110",
    "1111101111000001",
    "1111101101001101",
    "1111101101101110",
    "1111110000011010",
    "1111110101000000",
    "1111111011001111",
    "1111111101001000",
    "1111110100011110",
    "1111101011000000",
    "1111100001000011",
    "1111010110111100",
    "1111001101000101",
    "1111000011110110",
    "1110111011100101",
    "1110110100100100",
    "1110101111001000",
    "1110101011100101",
    "1110101010001011",
    "1110101011000111",
    "1110101110100001",
    "1110110100000101",
    "1110111011010100",
    "1111000011101010",
    "1111001100100001",
    "1111010101011111",
    "1111011110011111",
    "1111100111100101",
    "1111110000111000",
    "1111111010010100",
    "1111111100011100",
    "1111110100001000",
    "1111101101100101",
    "1111101001100101",
    "1111101000101000",
    "1111101010111010",
    "1111110000010100",
    "1111111000100111",
    "1111111100011110",
    "1111101111011010",
    "1111100000111001",
    "1111010010000011",
    "1111000100011000",
    "1110111001010110",
    "1110110010001011",
    "1110101111010111",
    "1110110000101011",
    "1110110101010010",
    "1110111100000101",
    "1111000100001011",
    "1111001100111101",
    "1111010110001001",
    "1111011111101100",
    "1111101001011001",
    "1111110010110010",
    "1111111011001001",
    "1111111110001010",
    "1111111001101001",
    "1111110111010000",
    "1111110110100010",
    "1111110110101101",
    "1111110110111100",
    "1111110110100111",
    "1111110101010110",
    "1111110011000110",
    "1111110000000000",
    "1111101100010111",
    "1111101000100010",
    "1111100100111110",
    "1111100010001000",
    "1111100000011010",
    "1111100000001101",
    "1111100001110011",
    "1111100101011010",
    "1111101011001101",
    "1111110011010100",
    "1111111101110001",
    "1111110101100000",
    "1111100110111101",
    "1111010111010101",
    "1111000111100111",
    "1110111001000001",
    "1110101100100101",
    "1110100011000000",
    "1110011100100110",
    "1110011001010001",
    "1110011000101000",
    "1110011010001110",
    "1110011101101101",
    "1110100010101111",
    "1110101001001011",
    "1110110000110101",
    "1110111001100011",
    "1111000011001011",
    "1111001101100110",
    "1111011000100010",
    "1111100011101010",
    "1111101110100000",
    "1111111000011010",
    "1111111111010111",
    "1111111001100101",
    "1111110110101100",
    "1111110110101010",
    "1111111000110111",
    "1111111100001001",
    "1111111111000001",
    "1111111111111110",
    "1111111101101111",
    "1111110111011101",
    "1111101100111110",
    "1111011110111111",
    "1111001110111010",
    "1110111110110101",
    "1110110001000010",
    "1110100111011000",
    "1110100011001101",
    "1110100100110110",
    "1110101011111010",
    "1110110111101010",
    "1111000111010011",
    "1111011010001100",
    "1111101111011100",
    "1111111010011000",
    "1111100101100010",
    "1111010100011000",
    "1111001000111111",
    "1111000100011000",
    "1111000110001000",
    "1111001100011100",
    "1111010100111011",
    "1111011101010100",
    "1111100100001101",
    "1111101001001111",
    "1111101100110111",
    "1111101111110101",
    "1111110010101011",
    "1111110101100101",
    "1111111000010100",
    "1111111010100010",
    "1111111011111010",
    "1111111100011001",
    "1111111100001000",
    "1111111011010111",
    "1111111010010000",
    "1111111000110111",
    "1111110111000110",
    "1111110100111101",
    "1111110010100011",
    "1111110000000101",
    "1111101101110000",
    "1111101011110001",
    "1111101010001011",
    "1111101000111000",
    "1111100111101011",
    "1111100110011110",
    "1111100101010010",
    "1111100100010011",
    "1111100011111110",
    "1111100100101001",
    "1111100110101110",
    "1111101010011011",
    "1111101111111001",
    "1111110111001100",
    "1111111111101010",
    "1111110100110011",
    "1111101000010100",
    "1111011010011110",
    "1111001011110010",
    "1110111101000000",
    "1110101111001100",
    "1110100011011100",
    "1110011010110000",
    "1110010101110001",
    "1110010100100101",
    "1110010110101010",
    "1110011010111010",
    "1110100000000011",
    "1110100100111001",
    "1110101000100000",
    "1110101010010110",
    "1110101010010001",
    "1110101000011011",
    "1110100101001101",
    "1110100001001101",
    "1110011101001111",
    "1110011010001001",
    "1110011000101010",
    "1110011001011001",
    "1110011100110101",
    "1110100011001000",
    "1110101100001111",
    "1110110111111001",
    "1111000101010101",
    "1111010011100010",
    "1111100001001100",
    "1111101100110111",
    "1111110101011000",
    "1111111001111101",
    "1111111010100000",
    "1111110111011100",
    "1111110001101001",
    "1111101010001001",
    "1111100001111011",
    "1111011001110111",
    "1111010010100100",
    "1111001100100001",
    "1111001000000100",
    "1111000101011101",
    "1111000100111011",
    "1111000110100010",
    "1111001010001100",
    "1111001111101011",
    "1111010110011101",
    "1111011101111111",
    "1111100101100010",
    "1111101100011100",
    "1111110010000110",
    "1111110110001000",
    "1111111000010100",
    "1111111000110011",
    "1111110111110110",
    "1111110101111001",
    "1111110011011001",
    "1111110000101111",
    "1111101110001110",
    "1111101100000110",
    "1111101010011110",
    "1111101001011001",
    "1111101000110111",
    "1111101000110101",
    "1111101001010010",
    "1111101010010000",
    "1111101011111100",
    "1111101110100000",
    "1111110010000110",
    "1111110110101001",
    "1111111011110001",
    "1111111111010001",
    "1111111011100001",
    "1111111001111011",
    "1111111011001101",
    "1111111111110001",
    "1111111000011110",
    "1111101110000100",
    "1111100001100100",
    "1111010011101110",
    "1111000101011101",
    "1110110111110111",
    "1110101100010100",
    "1110100100000110",
    "1110100000010111",
    "1110100001100110",
    "1110100111100101",
    "1110110001011111",
    "1110111101111000",
    "1111001011001111",
    "1111011000010101",
    "1111100100001010",
    "1111101110010101",
    "1111110110110111",
    "1111111110000100",
    "1111111011100001",
    "1111110101100001",
    "1111101111100001",
    "1111101001010111",
    "1111100011001010",
    "1111011101000100",
    "1111010111011011",
    "1111010010101001",
    "1111001110111011",
    "1111001100011110",
    "1111001011001110",
    "1111001011000111",
    "1111001100001111",
    "1111001110101001",
    "1111010010101100",
    "1111011000101101",
    "1111100001001000",
    "1111101100001100",
    "1111111001110100",
    "1111110110101011",
    "1111100110110001",
    "1111011000001110",
    "1111001100110011",
    "1111000101101111",
    "1111000011011000",
    "1111000101001001",
    "1111001001110101",
    "1111001111111011",
    "1111010110011000",
    "1111011100100110",
    "1111100010011100",
    "1111101000000000",
    "1111101101011011",
    "1111110010100010",
    "1111110110111101",
    "1111111010001100",
    "1111111011111001",
    "1111111011111110",
    "1111111010110110",
    "1111111001000111",
    "1111110111100111",
    "1111110111000100",
    "1111110111111101",
    "1111111010100101",
    "1111111110111101",
    "1111111011000010",
    "1111110011111001",
    "1111101100001010",
    "1111100100101010",
    "1111011110010111",
    "1111011010001110",
    "1111011001000100",
    "1111011011010110",
    "1111100001010000",
    "1111101010011100",
    "1111110110001110",
    "1111111100011100",
    "1111101110110111",
    "1111100010010000",
    "1111010111101100",
    "1111001111111011",
    "1111001011011001",
    "1111001010000111",
    "1111001011111100",
    "1111010000010111",
    "1111010110111011",
    "1111011111001100",
    "1111101000110010",
    "1111110011010111",
    "1111111110100111",
    "1111110101111000",
    "1111101010101110",
    "1111100000011110",
    "1111010111100111",
    "1111010000011111",
    "1111001011001010",
    "1111000111011010",
    "1111000100110011",
    "1111000010111011",
    "1111000001011010",
    "1111000000000111",
    "1110111110111111",
    "1110111110001001",
    "1110111101101011",
    "1110111101110010",
    "1110111110100001",
    "1110111111111010",
    "1111000001111110",
    "1111000100101110",
    "1111001000000110",
    "1111001100001110",
    "1111010001000010",
    "1111010110100101",
    "1111011100111100",
    "1111100100000000",
    "1111101011101101",
    "1111110011111010",
    "1111111100010100",
    "1111111011011101",
    "1111110100000000",
    "1111101101110101",
    "1111101001100001",
    "1111100111011101",
    "1111100111101110",
    "1111101010000010",
    "1111101101110001",
    "1111110010001010",
    "1111110110011011",
    "1111111010000000",
    "1111111101001011",
    "1111111110011101",
    "1111110110010010",
    "1111100111110111",
    "1111010010011001",
    "1110110111101101",
    "1110011100000100",
    "1110000100110001",
    "1101110110100000",
    "1101110011010111",
    "1101111010001111",
    "1110000111011010",
    "1110010110001000",
    "1110100010100010",
    "1110101010101010",
    "1110101110011100",
    "1110101111010100",
    "1110101111000111",
    "1110101111001010",
    "1110110000001000",
    "1110110010000110",
    "1110110100110111",
    "1110111000011000",
    "1110111100110101",
    "1111000010100010",
    "1111001001011110",
    "1111010001010000",
    "1111011001001100",
    "1111100000100110",
    "1111100111000100",
    "1111101100010101",
    "1111110000010011",
    "1111110010111111",
    "1111110100011101",
    "1111110100111111",
    "1111110100111110",
    "1111110100110011",
    "1111110100110100",
    "1111110101000111",
    "1111110101011010",
    "1111110100111011",
    "1111110010101100",
    "1111101101101011",
    "1111100101001011",
    "1111011001001100",
    "1111001010101011",
    "1110111011011000",
    "1110101101011011",
    "1110100010101011",
    "1110011100001001",
    "1110011001111010",
    "1110011011001001",
    "1110011110101000",
    "1110100011010000",
    "1110101000001110",
    "1110101101001010",
    "1110110010001011",
    "1110110111101101",
    "1110111110001100",
    "1111000110000001",
    "1111001111011001",
    "1111011010001111",
    "1111100110001101",
    "1111110010011000",
    "1111111101100000",
    "1111111001110111",
    "1111110101001101",
    "1111110101011010",
    "1111111010100011",
    "1111111100001111",
    "1111110000110101",
    "1111100101100010",
    "1111011100101010",
    "1111010111111111",
    "1111011000011101",
    "1111011110000010",
    "1111101000000101",
    "1111110101010110",
    "1111111011100011",
    "1111101100000000",
    "1111011101001010",
    "1111001111111011",
    "1111000101000101",
    "1110111101000000",
    "1110110111111010",
    "1110110101101010",
    "1110110101110110",
    "1110110111110001",
    "1110111010101011",
    "1110111101111010",
    "1111000000111001",
    "1111000011010101",
    "1111000101000110",
    "1111000110001011",
    "1111000110011111",
    "1111000101111110",
    "1111000100100000",
    "1111000010000011",
    "1110111110101110",
    "1110111010111010",
    "1110110111001001",
    "1110110100001110",
    "1110110010110110",
    "1110110011100111",
    "1110110110110100",
    "1110111100011011",
    "1111000100000001",
    "1111001101000111",
    "1111010111001000",
    "1111100001100111",
    "1111101100011101",
    "1111110111100111",
    "1111111100111001",
    "1111110001011000",
    "1111100110011010",
    "1111011100110111",
    "1111010101100111",
    "1111010001010101",
    "1111010000001101",
    "1111010001110100",
    "1111010101011010",
    "1111011010000100",
    "1111011111000101",
    "1111100100001101",
    "1111101001100101",
    "1111101111101100",
    "1111110111000101",
    "1111111111111001",
    "1111110101011010",
    "1111101010001000",
    "1111011111010010",
    "1111010110100100",
    "1111010001100001",
    "1111010001011100",
    "1111010110101100",
    "1111100000100001",
    "1111101101001101",
    "1111111010010011",
    "1111111010101011",
    "1111110011111000",
    "1111110010011010",
    "1111110110100001",
    "1111111111100011",
    "1111110011101010",
    "1111100100110111",
    "1111010101111001",
    "1111001000100010",
    "1110111110010110",
    "1110111000010000",
    "1110110110100100",
    "1110111000110101",
    "1110111110001101",
    "1111000101100100",
    "1111001101110010",
    "1111010110001011",
    "1111011110010110",
    "1111100110000011",
    "1111101101000110",
    "1111110011010010",
    "1111111000011000",
    "1111111100000111",
    "1111111110011010",
    "1111111111010101",
    "1111111111000110",
    "1111111110001011",
    "1111111100111100",
    "1111111011110011",
    "1111111011000011",
    "1111111010111010",
    "1111111011100100",
    "1111111101001001",
    "1111111111101111",
    "1111111100100011",
    "1111110111110101",
    "1111110010000110",
    "1111101011100011",
    "1111100100011010",
    "1111011101000111",
    "1111010110001001",
    "1111010000000111",
    "1111001011011110",
    "1111001000101010",
    "1111000111111001",
    "1111001001001001",
    "1111001100010001",
    "1111010001000010",
    "1111010111001110",
    "1111011110101101",
    "1111100111011110",
    "1111110001101001",
    "1111111101010101",
    "1111110101100000",
    "1111100111010100",
    "1111011000110100",
    "1111001011000001",
    "1110111111000010",
    "1110110101110010",
    "1110101111111011",
    "1110101101101001",
    "1110101110110101",
    "1110110011001101",
    "1110111010010011",
    "1111000011101001",
    "1111001110011110",
    "1111011001110101",
    "1111100100100010",
    "1111101101010100",
    "1111110011010011",
    "1111110110000111",
    "1111110110000000",
    "1111110011101111",
    "1111110000010001",
    "1111101100010101",
    "1111101000001010",
    "1111100011011111",
    "1111011101101001",
    "1111010110010000",
    "1111001101011110",
    "1111000100001101",
    "1110111011110011",
    "1110110101100101",
    "1110110010100001",
    "1110110010101110",
    "1110110101100100",
    "1110111010000100",
    "1110111111000101",
    "1111000011111000",
    "1111001000000001",
    "1111001011100001",
    "1111001110011011",
    "1111010000110011",
    "1111010010100111",
    "1111010011101110",
    "1111010100000011",
    "1111010011101001",
    "1111010010101001",
    "1111010001010101",
    "1111010000000010",
    "1111001111000000",
    "1111001110100001",
    "1111001110111000",
    "1111010000011001",
    "1111010011010011",
    "1111010111110100",
    "1111011101111010",
    "1111100101011000",
    "1111101101110100",
    "1111110110110000",
    "1111111111101010",
    "1111110111111101",
    "1111110000101001",
    "1111101010110101",
    "1111100110110111",
    "1111100100111110",
    "1111100101011000",
    "1111101000001010",
    "1111101101010100",
    "1111110100110011",
    "1111111110010110",
    "1111110110011111",
    "1111101010101111",
    "1111011111101000",
    "1111010110101000",
    "1111010001010100",
    "1111010000111110",
    "1111010110011111",
    "1111100001111110",
    "1111110010101011",
    "1111111001001101",
    "1111100100010000",
    "1111010001001000",
    "1111000010000101",
    "1110111000011000",
    "1110110100000110",
    "1110110100011010",
    "1110110111111010",
    "1110111101011011",
    "1111000100001010",
    "1111001011111010",
    "1111010100101010",
    "1111011110010001",
    "1111101000000000",
    "1111110000110001",
    "1111110111000100",
    "1111111001100101",
    "1111110111110001",
    "1111110001111111",
    "1111101001101000",
    "1111100000100110",
    "1111011000111100",
    "1111010100010000",
    "1111010011100001",
    "1111010110110111",
    "1111011110000000",
    "1111101000001000",
    "1111110100000111",
    "1111111111000111",
    "1111110010110111",
    "1111101000001010",
    "1111011111110110",
    "1111011010011110",
    "1111011000000100",
    "1111011000011000",
    "1111011010110101",
    "1111011110110011",
    "1111100011101111",
    "1111101001011011",
    "1111101111110100",
    "1111110111000011",
    "1111111111010011",
    "1111110111010011",
    "1111101100111111",
    "1111100010000000",
    "1111010110110111",
    "1111001100001110",
    "1111000010101110",
    "1110111011000010",
    "1110110101011101",
    "1110110010000011",
    "1110110000100011",
    "1110110000011110",
    "1110110001010101",
    "1110110010111001",
    "1110110101001011",
    "1110111000011110",
    "1110111101011001",
    "1111000100110110",
    "1111001111111111",
    "1111011111101110",
    "1111110100000011",
    "1111110100011010",
    "1111011100011011",
    "1111000111001101",
    "1110110111100010",
    "1110101110111000",
    "1110101101001001",
    "1110110000110101",
    "1110110111111100",
    "1111000001001000",
    "1111001011111111",
    "1111011000110000",
    "1111100111100000",
    "1111110111010100",
    "1111111001110001",
    "1111101110010100",
    "1111101000100001",
    "1111101001001011",
    "1111101111001110",
    "1111110111111001",
    "1111111111100111",
    "1111111100110011",
    "1111111111001110",
    "1111111000011011",
    "1111101011111010",
    "1111011101110000",
    "1111010000100100",
    "1111000110010010",
    "1110111111110110",
    "1110111101010001",
    "1110111101111011",
    "1111000001001111",
    "1111000110111011",
    "1111001111001111",
    "1111011010101010",
    "1111101001011110",
    "1111111011011100",
    "1111110000011111",
    "1111011100000101",
    "1111001001010001",
    "1110111001101000",
    "1110101110000101",
    "1110100110110001",
    "1110100011001101",
    "1110100010110100",
    "1110100101001101",
    "1110101010010001",
    "1110110010001010",
    "1110111100110000",
    "1111001001011101",
    "1111010111000001",
    "1111100011111001",
    "1111101110100101",
    "1111110110001100",
    "1111111010101110",
    "1111111101000101",
    "1111111110110010",
    "1111111110010110",
    "1111111000110100",
    "1111101111100100",
    "1111100010100100",
    "1111010010111101",
    "1111000010111011",
    "1110110101001000",
    "1110101100000001",
    "1110101001001100",
    "1110101101000100",
    "1110110110101010",
    "1111000011111000",
    "1111010010001101",
    "1111011111001111",
    "1111101001000110",
    "1111101110111000",
    "1111110000110100",
    "1111110000001111",
    "1111101111001011",
    "1111101111110100",
    "1111110011111010",
    "1111111100010101",
    "1111110111000100",
    "1111100111101010",
    "1111010111100000",
    "1111001001000001",
    "1110111110010111",
    "1110111000111110",
    "1110111001001110",
    "1110111110011011",
    "1111000110111110",
    "1111010001000000",
    "1111011010110010",
    "1111100011000110",
    "1111101001100000",
    "1111101110010001",
    "1111110010001100",
    "1111110110010110",
    "1111111011110100",
    "1111111100011110",
    "1111110010000000",
    "1111100100101111",
    "1111010101011010",
    "1111000101100000",
    "1110110111001011",
    "1110101100100110",
    "1110100111100101",
    "1110101001001011",
    "1110110001001111",
    "1110111110101110",
    "1111001111111010",
    "1111100010101100",
    "1111110101000011",
    "1111111010110010",
    "1111101110001101",
    "1111100101111100",
    "1111100001111110",
    "1111100001100111",
    "1111100011100111",
    "1111100110101001",
    "1111101001101110",
    "1111101100011111",
    "1111101111010011",
    "1111110011000001",
    "1111111000110000",
    "1111111110100000",
    "1111110010010010",
    "1111100010011010",
    "1111001111011001",
    "1110111010100101",
    "1110100110000001",
    "1110010100010010",
    "1110000111110100",
    "1110000010001101",
    "1110000011110110",
    "1110001011101101",
    "1110010111100101",
    "1110100100111011",
    "1110110001100110",
    "1110111100001001",
    "1111000100000110",
    "1111001001011110",
    "1111001100101101",
    "1111001110001100",
    "1111001110011111",
    "1111001110001101",
    "1111001110000101",
    "1111001110111000",
    "1111010001010000",
    "1111010101100101",
    "1111011011111000",
    "1111100011101111",
    "1111101100100101",
    "1111110101111001",
    "1111111111010110",
    "1111110111010000",
    "1111101110000101",
    "1111100101001101",
    "1111011100101011",
    "1111010100100100",
    "1111001101000000",
    "1111000110001001",
    "1111000000011001",
    "1110111100001110",
    "1110111010010011",
    "1110111011001010",
    "1110111111010001",
    "1111000110101010",
    "1111010001000000",
    "1111011101110010",
    "1111101100001101",
    "1111111011100110",
    "1111110100101110",
    "1111100101011111",
    "1111010111011011",
    "1111001011011011",
    "1111000010010100",
    "1110111100110010",
    "1110111011000100",
    "1110111100101011",
    "1111000000011111",
    "1111000101000001",
    "1111001000101111",
    "1111001010101011",
    "1111001010100011",
    "1111001000101000",
    "1111000101110001",
    "1111000010111001",
    "1111000000110011",
    "1110111111111010",
    "1111000000001101",
    "1111000001010101",
    "1111000010101011",
    "1111000011100001",
    "1111000011011000",
    "1111000010000010",
    "1110111111100100",
    "1110111100100101",
    "1110111001111111",
    "1110111001010101",
    "1110111100010001",
    "1111000100001000",
    "1111010001001000",
    "1111100010001000",
    "1111110100111101",
    "1111111001001011",
    "1111101011000100",
    "1111100010101001",
    "1111100000100100",
    "1111100100011000",
    "1111101100110001",
    "1111111000000011",
    "1111111011011011",
    "1111101111011000",
    "1111100101010000",
    "1111011110010010",
    "1111011011011000",
    "1111011100111000",
    "1111100010100111",
    "1111101011110100",
    "1111110111001101",
    "1111111100100100",
    "1111110000101111",
    "1111100101110110",
    "1111011100000010",
    "1111010011000011",
    "1111001010101101",
    "1111000011000011",
    "1110111100011001",
    "1110110111001011",
    "1110110011111001",
    "1110110010111001",
    "1110110100010011",
    "1110110111111111",
    "1110111101101000",
    "1111000100100101",
    "1111001100001010",
    "1111010011011100",
    "1111011001100010",
    "1111011101100110",
    "1111011111010010",
    "1111011110110011",
    "1111011100111000",
    "1111011010111000",
    "1111011010001100",
    "1111011100000100",
    "1111100001000111",
    "1111101001001100",
    "1111110011011101",
    "1111111110101010",
    "1111110110100010",
    "1111101101011001",
    "1111100110110001",
    "1111100011001000",
    "1111100010100110",
    "1111100100111110",
    "1111101001110100",
    "1111110000100011",
    "1111111000011101",
    "1111111111001001",
    "1111110111000011",
    "1111101111101010",
    "1111101001001111",
    "1111100011101010",
    "1111011110100011",
    "1111011001001100",
    "1111010010100001",
    "1111001001001011",
    "1110111011111101",
    "1110101010100110",
    "1110010110010011",
    "1110000001100001",
    "1101101111010100",
    "1101100010100110",
    "1101011101000010",
    "1101011110110000",
    "1101100110001001",
    "1101110000110101",
    "1101111100101010",
    "1110001000110101",
    "1110010110000011",
    "1110100101101111",
    "1110111000111100",
    "1111001111010110",
    "1111100110111110",
    "1111111100110000",
    "1111110010100100",
    "1111101001010000",
    "1111100111100111",
    "1111101100000011",
    "1111110011111001",
    "1111111100011100",
    "1111111100010100",
    "1111110111100000",
    "1111110101001110",
    "1111110100111110",
    "1111110101111111",
    "1111110111100010",
    "1111111001000110",
    "1111111010010010",
    "1111111010110000",
    "1111111010000011",
    "1111110111101110",
    "1111110011011101",
    "1111101101000001",
    "1111100100011010",
    "1111011001101000",
    "1111001100111100",
    "1110111111000101",
    "1110110001010111",
    "1110100101011011",
    "1110011100110010",
    "1110011000011010",
    "1110011000010001",
    "1110011011100011",
    "1110100000110110",
    "1110100110110010",
    "1110101100110000",
    "1110110010111101",
    "1110111010010001",
    "1111000011111001",
    "1111010000111001",
    "1111100001101001",
    "1111110101101110",
    "1111110100011000",
    "1111011110111111",
    "1111001100100000",
    "1110111110111000",
    "1110110111010001",
    "1110110101110001",
    "1110111001101000",
    "1111000001110001",
    "1111001101001100",
    "1111011011010100",
    "1111101100001111",
    "1111111111101101",
    "1111101000110101",
    "1111010000100001",
    "1110111001010101",
    "1110100110010010",
    "1110011001110111",
    "1110010101001101",
    "1110010111101000",
    "1110011111000100",
    "1110101000100111",
    "1110110001110011",
    "1110111001001011",
    "1110111110010111",
    "1111000001110000",
    "1111000011110011",
    "1111000100111001",
    "1111000101010101",
    "1111000101001101",
    "1111000100111011",
    "1111000101001011",
    "1111000110111110",
    "1111001011001111",
    "1111010010100111",
    "1111011100111101",
    "1111101001100001",
    "1111110111001111",
    "1111111010111100",
    "1111101101111010",
    "1111100010010000",
    "1111011000011011",
    "1111010000110001",
    "1111001011100110",
    "1111001001010000",
    "1111001001111001",
    "1111001101100000",
    "1111010011110011",
    "1111011100010100",
    "1111100110100101",
    "1111110010000100",
    "1111111110010011",
    "1111110101001001",
    "1111101000111101",
    "1111011101110010",
    "1111010100011000",
    "1111001101011011",
    "1111001001010001",
    "1111000111111110",
    "1111001001001100",
    "1111001100100001",
    "1111010001100001",
    "1111010111111110",
    "1111011111101100",
    "1111101000100111",
    "1111110010101001",
    "1111111101100011",
    "1111110110110110",
    "1111101010110100",
    "1111011110010111",
    "1111010001010111",
    "1111000011100111",
    "1110110101001000",
    "1110100110010011",
    "1110010111111110",
    "1110001011001111",
    "1110000001001111",
    "1101111010100101",
    "1101110111011000",
    "1101110111000011",
    "1101111000110111",
    "1101111100001010",
    "1110000000111001",
    "1110000111011111",
    "1110010000101001",
    "1110011101000000",
    "1110101100100001",
    "1110111110001111",
    "1111010000011010",
    "1111100000111110",
    "1111101110001010",
    "1111110110111010",
    "1111111011010010",
    "1111111100001110",
    "1111111011001001",
    "1111111001100110",
    "1111111000110101",
    "1111111001110001",
    "1111111100101101",
    "1111111110011100",
    "1111111000011001",
    "1111110010000001",
    "1111101100010011",
    "1111101000000111",
    "1111100110000110",
    "1111100110100101",
    "1111101001101010",
    "1111101111011110",
    "1111111000010011",
    "1111111011010010",
    "1111101010110000",
    "1111010101111001",
    "1110111101100001",
    "1110100011111011",
    "1110001100010110",
    "1101111010001100",
    "1101101111111111",
    "1101101110011110",
    "1101110100101001",
    "1110000000000000",
    "1110001101100110",
    "1110011010111101",
    "1110100110101000",
    "1110110000010010",
    "1110111000001011",
    "1110111110110110",
    "1111000100101001",
    "1111001001100011",
    "1111001101011001",
    "1111010000000010",
    "1111010001101001",
    "1111010010101111",
    "1111010100000101",
    "1111010110001110",
    "1111011001100000",
    "1111011101101001",
    "1111100010000110",
    "1111100110001001",
    "1111101001000101",
    "1111101010011001",
    "1111101001110010",
    "1111100111001011",
    "1111100010101001",
    "1111011100011110",
    "1111010101001000",
    "1111001101001111",
    "1111000101100100",
    "1110111110110011",
    "1110111001010101",
    "1110110101001001",
    "1110110001111110",
    "1110101111001010",
    "1110101100001110",
    "1110101000111100",
    "1110100101100111",
    "1110100010110110",
    "1110100001011010",
    "1110100010000000",
    "1110100100111100",
    "1110101010011101",
    "1110110010100010",
    "1110111101011011",
    "1111001011100000",
    "1111011101001111",
    "1111110010111100",
    "1111110100000011",
    "1111011001101010",
    "1111000000101100",
    "1110101100010011",
    "1110011110110101",
    "1110011001001110",
    "1110011010100110",
    "1110100000111001",
    "1110101001101000",
    "1110110010110011",
    "1110111011101000",
    "1111000100010010",
    "1111001101100001",
    "1111010111110001",
    "1111100010101011",
    "1111101101001011",
    "1111110101111010",
    "1111111011110000",
    "1111111110011110",
    "1111111110110011",
    "1111111110010010",
    "1111111110100101",
    "1111111111001001",
    "1111111010100010",
    "1111110100000000",
    "1111101100011111",
    "1111100101000011",
    "1111011110101101",
    "1111011010000100",
    "1111010111101000",
    "1111010111101010",
    "1111011010001110",
    "1111011111010010",
    "1111100110100101",
    "1111101111100011",
    "1111111001011010",
    "1111111100110000",
    "1111110011111110",
    "1111101101001000",
    "1111101000110011",
    "1111100111010010",
    "1111101000011011",
    "1111101011101001",
    "1111110000001000",
    "1111110100111111",
    "1111111001010111",
    "1111111100100000",
    "1111111101101110",
    "1111111100010111",
    "1111110111110011",
    "1111101111101011",
    "1111100100001011",
    "1111010110010101",
    "1111000111111001",
    "1110111011001111",
    "1110110010100111",
    "1110101111101001",
    "1110110011000000",
    "1110111100001111",
    "1111001010001100",
    "1111011011001010",
    "1111101101010000",
    "1111111110100101",
    "1111110010011111",
    "1111100111011010",
    "1111100001001111",
    "1111100000010111",
    "1111100100101111",
    "1111101101110110",
    "1111111011000011",
    "1111110100000011",
    "1111100000001010",
    "1111001010011101",
    "1110110100110110",
    "1110100001111000",
    "1110010100000000",
    "1110001100111111",
    "1110001101010110",
    "1110010100000110",
    "1110011111001010",
    "1110101100010001",
    "1110111001110111",
    "1111000111001011",
    "1111010100001000",
    "1111100000100110",
    "1111101011111110",
    "1111110101000101",
    "1111111010011001",
    "1111111010110010",
    "1111110110010000",
    "1111101110001101",
    "1111100101011000",
    "1111011111000000",
    "1111011101111000",
    "1111100011100100",
    "1111101111110100",
    "1111111111001011",
    "1111101100011101",
    "1111011011000001",
    "1111001101001010",
    "1111000011111001",
    "1110111110110011",
    "1110111100101011",
    "1110111100001111",
    "1110111100110011",
    "1110111110110011",
    "1111000011011000",
    "1111001100001010",
    "1111011010001111",
    "1111101101100011",
    "1111111011100000",
    "1111100011111001",
    "1111001110111000",
    "1110111111001010",
    "1110110110001000",
    "1110110011011111",
    "1110110101101100",
    "1110111010110000",
    "1111000001000101",
    "1111001000000001",
    "1111001111110011",
    "1111011000111111",
    "1111100011101100",
    "1111101110111101",
    "1111111000110100",
    "1111111110110000",
    "1111111110110000",
    "1111111000010000",
    "1111101100100000",
    "1111011110011110",
    "1111010001110100",
    "1111001001110111",
    "1111001000100011",
    "1111001110000111",
    "1111011001010001",
    "1111100111110110",
    "1111110111100011",
    "1111111001011100",
    "1111101100010100",
    "1111100001011010",
    "1111011000110000",
    "1111010010010000",
    "1111001110001001",
    "1111001100111000",
    "1111001111001101",
    "1111010101101001",
    "1111100000001100",
    "1111101101111001",
    "1111111100111010",
    "1111110101011010",
    "1111101011110001",
    "1111101000000101",
    "1111101010111101",
    "1111110011011111",
    "1111111111100111",
    "1111110011001001",
    "1111100111000001",
    "1111011101001111",
    "1111010110001000",
    "1111010001100001",
    "1111001111001111",
    "1111001111100001",
    "1111010011000001",
    "1111011010100010",
    "1111100110001110",
    "1111110101010111",
    "1111111001111101",
    "1111101010011011",
    "1111011110101011",
    "1111011000100101",
    "1111011000110100",
    "1111011110111010",
    "1111101001011101",
    "1111110110110100",
    "1111111010101001",
    "1111101100100011",
    "1111100000010010",
    "1111010111010011",
    "1111010011000001",
    "1111010100101001",
    "1111011100111111",
    "1111101100000000",
    "1111111111001101",
    "1111100110110000",
    "1111001101010100",
    "1110110101110010",
    "1110100010101011",
    "1110010101100000",
    "1110001110110011",
    "1110001110000101",
    "1110010010011111",
    "1110011011001010",
    "1110100111101010",
    "1110110111111001",
    "1111001011101000",
    "1111100010000010",
    "1111111001001001",
    "1111110001110010",
    "1111100001111001",
    "1111011001011110",
    "1111011001011000",
    "1111100000101001",
    "1111101100110011",
    "1111111010100111",
    "1111111000111100",
    "1111110000001101",
    "1111101100001101",
    "1111101100111100",
    "1111110001100110",
    "1111111001000011",
    "1111111101101111",
    "1111110011101001",
    "1111101001000011",
    "1111011110001111",
    "1111010011011111",
    "1111001001011001",
    "1111000000111001",
    "1110111011001001",
    "1110111001010001",
    "1110111100001001",
    "1111000100000011",
    "1111010000011110",
    "1111100000001000",
    "1111110001011001",
    "1111111101011110",
    "1111101101111001",
    "1111100000011010",
    "1111010100111110",
    "1111001011001010",
    "1111000010101001",
    "1110111011011110",
    "1110110110000100",
    "1110110011000011",
    "1110110010111000",
    "1110110101011111",
    "1110111010011000",
    "1111000000101001",
    "1111000111100011",
    "1111001110111010",
    "1111010111010000",
    "1111100001101001",
    "1111101111000100",
    "1111111111011001",
    "1111101110110100",
    "1111011110001101",
    "1111010001011111",
    "1111001010101010",
    "1111001010010110",
    "1111001111111010",
    "1111011001110101",
    "1111100110101000",
    "1111110100111101",
    "1111111100010101",
    "1111101110110011",
    "1111100100001011",
    "1111011110011100",
    "1111011111001101",
    "1111100111010100",
    "1111110101111001",
    "1111110111010110",
    "1111100011111100",
    "1111010011011111",
    "1111001000101101",
    "1111000100111001",
    "1111000111111010",
    "1111010000100110",
    "1111011101110010",
    "1111101110110011",
    "1111111100110001",
    "1111100101111001",
    "1111001110010110",
    "1110111000100101",
    "1110100111001011",
    "1110011100000010",
    "1110010111110001",
    "1110011001101011",
    "1110100000001101",
    "1110101001101101",
    "1110110101001001",
    "1111000010010111",
    "1111010001110001",
    "1111100011101010",
    "1111110111101100",
    "1111110011100110",
    "1111100000100110",
    "1111010001111000",
    "1111001001100000",
    "1111001000011101",
    "1111001110011111",
    "1111011010001100",
    "1111101001100010",
    "1111111010001110",
    "1111110101111111",
    "1111101001010000",
    "1111100001001010",
    "1111011110011011",
    "1111100000110101",
    "1111100111010101",
    "1111110000100101",
    "1111111011001101",
    "1111111001110100",
    "1111101111100000",
    "1111100110111000",
    "1111100001001100",
    "1111011111101110",
    "1111100011011010",
    "1111101100011000",
    "1111111001101000",
    "1111110110111000",
    "1111100111110110",
    "1111011011110000",
    "1111010100010010",
    "1111010001111001",
    "1111010100000001",
    "1111011001011101",
    "1111100001001000",
    "1111101010011001",
    "1111110100111111",
    "1111111111001101",
    "1111110011000011",
    "1111101000000010",
    "1111100000010010",
    "1111011101100110",
    "1111100000110101",
    "1111101001001101",
    "1111110100110100",
    "1111111111000001",
    "1111110100110110",
    "1111101110001111",
    "1111101011101101",
    "1111101100110101",
    "1111110000111000",
    "1111110111001010",
    "1111111111010001",
    "1111110111000000",
    "1111101100010111",
    "1111100010001000",
    "1111011010011000",
    "1111010111011000",
    "1111011010110111",
    "1111100101000101",
    "1111110100101101",
    "1111111000101110",
    "1111100110010101",
    "1111010110101100",
    "1111001011010100",
    "1111000100101110",
    "1111000010101001",
    "1111000100100101",
    "1111001010000100",
    "1111010010101111",
    "1111011110010010",
    "1111101100000111",
    "1111111011010001",
    "1111110101100011",
    "1111100111111111",
    "1111011101100001",
    "1111010111001001",
    "1111010101001101",
    "1111010111001001",
    "1111011011111000",
    "1111100001111011",
    "1111100111011100",
    "1111101010101110",
    "1111101010010010",
    "1111100101010011",
    "1111011011101111",
    "1111001110100001",
    "1110111111010111",
    "1110110000010111",
    "1110100011010111",
    "1110011001100101",
    "1110010011010010",
    "1110010000000111",
    "1110001111010110",
    "1110010000011100",
    "1110010011001111",
    "1110010111111111",
    "1110011111010010",
    "1110101001100011",
    "1110110110101010",
    "1111000101110010",
    "1111010101100000",
    "1111100100000101",
    "1111101111101110",
    "1111110111000011",
    "1111111001000101",
    "1111110101011010",
    "1111101100001101",
    "1111011110011100",
    "1111001101110000",
    "1110111100011001",
    "1110101100101110",
    "1110100001000000",
    "1110011010111000",
    "1110011011011011",
    "1110100010111011",
    "1110110001000010",
    "1111000100011010",
    "1111011010111010",
    "1111110001100111",
    "1111111010100001",
    "1111101100001000",
    "1111100100110110",
    "1111100101000001",
    "1111101011111110",
    "1111111000000111",
    "1111111000110000",
    "1111101001010100",
    "1111011100000111",
    "1111010011011101",
    "1111010000110101",
    "1111010100101111",
    "1111011110100011",
    "1111101100100111",
    "1111111100101010",
    "1111110011011101",
    "1111100101101110",
    "1111011011010001",
    "1111010100111011",
    "1111010011001000",
    "1111010110010101",
    "1111011110110001",
    "1111101100010000",
    "1111111101101001",
    "1111101111000111",
    "1111011100110000",
    "1111001101101011",
    "1111000011011010",
    "1110111110001101",
    "1110111101010100",
    "1110111111010001",
    "1111000010101110",
    "1111000110110001",
    "1111001011000001",
    "1111001111010110",
    "1111010011011010",
    "1111010110011101",
    "1111010111011000",
    "1111010101001000",
    "1111001111001000",
    "1111000101100100",
    "1110111001011001",
    "1110101100010111",
    "1110100000010101",
    "1110010110111110",
    "1110010001100010",
    "1110010000110110",
    "1110010101011101",
    "1110011111110000",
    "1110101111110001",
    "1111000101000011",
    "1111011110010010",
    "1111111001011110",
    "1111101100000011",
    "1111010101001001",
    "1111000100010101",
    "1110111011010001",
    "1110111010101011",
    "1111000010001010",
    "1111010000010010",
    "1111100010111000",
    "1111110111010000",
    "1111110101010010",
    "1111100101001110",
    "1111011010000111",
    "1111010100100111",
    "1111010100011101",
    "1111011001001001",
    "1111100010011001",
    "1111110000010110",
    "1111111100110111",
    "1111100110001110",
    "1111001101111101",
    "1110110111100011",
    "1110100111000011",
    "1110011111111010",
    "1110100100001101",
    "1110110011101001",
    "1111001011011011",
    "1111100111001000",
    "1111111110000110",
    "1111101000010001",
    "1111011001100011",
    "1111010010010101",
    "1111010001011100",
    "1111010101000000",
    "1111011011010100",
    "1111100011011000",
    "1111101100110010",
    "1111110111011001",
    "1111111100110110",
    "1111110000011011",
    "1111100100000001",
    "1111011000101100",
    "1111001111011110",
    "1111001001010001",
    "1111000110100100",
    "1111000110111110",
    "1111001001101010",
    "1111001101100011",
    "1111010001110000",
    "1111010101100111",
    "1111011000111010",
    "1111011011101111",
    "1111011110001100",
    "1111100000011111",
    "1111100010100111",
    "1111100100001101",
    "1111100100101001",
    "1111100011001111",
    "1111011111101100",
    "1111011010011000",
    "1111010100001110",
    "1111001110101110",
    "1111001011001111",
    "1111001010101011",
    "1111001100111100",
    "1111010001001000",
    "1111010101110010",
    "1111011001100010",
    "1111011011010011",
    "1111011010101111",
    "1111011000001100",
    "1111010100100100",
    "1111010000111000",
    "1111001101111011",
    "1111001100001001",
    "1111001011100000",
    "1111001011101111",
    "1111001100011100",
    "1111001100111010",
    "1111001100001111",
    "1111001001011011",
    "1111000011100100",
    "1110111010011001",
    "1110101110010111",
    "1110100000110000",
    "1110010011011100",
    "1110001000011101",
    "1110000001001111",
    "1101111110011011",
    "1101111111101001",
    "1110000011111110",
    "1110001010001100",
    "1110010001100100",
    "1110011010000110",
    "1110100100010101",
    "1110110001000101",
    "1111000000101001",
    "1111010010011010",
    "1111100100110111",
    "1111110110000101",
    "1111111011100111",
    "1111110001010010",
    "1111101010111001",
    "1111100111101110",
    "1111100110111001",
    "1111100111111101",
    "1111101011010011",
    "1111110010000111",
    "1111111101110010",
    "1111110001001000",
    "1111011011110011",
    "1111000101000110",
    "1110110001000011",
    "1110100011110001",
    "1110100000000011",
    "1110100110101000",
    "1110110101110001",
    "1111001010001001",
    "1111011111110011",
    "1111110011011100",
    "1111111100111101",
    "1111110010001000",
    "1111101011101101",
    "1111101000111001",
    "1111101001000011",
    "1111101011110100",
    "1111110001001000",
    "1111111000110000",
    "1111111101110100",
    "1111110011110101",
    "1111101010110010",
    "1111100100001101",
    "1111100001001100",
    "1111100010001000",
    "1111100110101110",
    "1111101110001100",
    "1111110111100011",
    "1111111110000101",
    "1111110011011101",
    "1111101000111000",
    "1111011110101000",
    "1111010101001011",
    "1111001101010111",
    "1111001000011000",
    "1111000111011011",
    "1111001011010100",
    "1111010100001101",
    "1111100001000111",
    "1111110000010011",
    "1111111111101110",
    "1111110010011001",
    "1111100111001110",
    "1111011110110011",
    "1111011000010001",
    "1111010010011101",
    "1111001100011100",
    "1111000110001001",
    "1111000000010100",
    "1110111100000100",
    "1110111010011000",
    "1110111011011101",
    "1110111110011111",
    "1111000010001011",
    "1111000101001011",
    "1111000110110100",
    "1111000111011111",
    "1111001000100000",
    "1111001011100000",
    "1111010001110100",
    "1111011011101101",
    "1111101000010000",
    "1111110101100011",
    "1111111110100110",
    "1111110101111111",
    "1111110001001011",
    "1111101111100000",
    "1111101111100000",
    "1111101111110000",
    "1111101111101011",
    "1111101111110010",
    "1111110001010010",
    "1111110101011001",
    "1111111100100010",
    "1111111010000111",
    "1111110000101110",
    "1111101001110000",
    "1111100111010010",
    "1111101010000110",
    "1111110001011000",
    "1111111010111101",
    "1111111011110000",
    "1111110101000000",
    "1111110001110000",
    "1111110001100100",
    "1111110011000111",
    "1111110101000000",
    "1111110110101101",
    "1111111000101101",
    "1111111100001011",
    "1111111101110110",
    "1111110101100001",
    "1111101100010000",
    "1111100100111110",
    "1111100011001111",
    "1111101010001010",
    "1111111011000010",
    "1111101011100110",
    "1111001101110010",
    "1110110000110000",
    "1110011001010110",
    "1110001010100000",
    "1110000100100101",
    "1110000101101010",
    "1110001010110000",
    "1110010001100001",
    "1110011001011101",
    "1110100100001011",
    "1110110100000000",
    "1111001010000111",
    "1111100101010011",
    "1111111110001010",
    "1111100101011101",
    "1111010101001101",
    "1111001111110110",
    "1111010100100100",
    "1111011111101000",
    "1111101011110011",
    "1111110100101000",
    "1111110111101101",
    "1111110101010100",
    "1111101111101011",
    "1111101001110101",
    "1111100110010101",
    "1111100110010011",
    "1111101001000011",
    "1111101100101101",
    "1111101111001000",
    "1111101111000000",
    "1111101100100001",
    "1111101001011111",
    "1111101000111100",
    "1111101110010010",
    "1111111100000000",
    "1111101101100101",
    "1111010001001010",
    "1110110011100111",
    "1110011010100010",
    "1110001010000110",
    "1110000011100010",
    "1110000100110100",
    "1110001001100010",
    "1110001101000101",
    "1110001100101110",
    "1110001000100101",
    "1110000011100010",
    "1110000001100111",
    "1110000110000011",
    "1110010001010101",
    "1110100000110011",
    "1110101111100011",
    "1110111000100111",
    "1110111001000110",
    "1110110001011100",
    "1110100101011000",
    "1110011010100000",
    "1110010110010010",
    "1110011011110011",
    "1110101010111010",
    "1111000000010101",
    "1111010111000100",
    "1111101010001010",
    "1111110110011011",
    "1111111011100100",
    "1111111011111110",
    "1111111011011010",
    "1111111101000001",
    "1111111110000101",
    "1111110111101010",
    "1111110011100100",
    "1111110110000101",
    "1111111110001101",
    "1111101010000110",
    "1111010001010111",
    "1110111001101011",
    "1110101000101000",
    "1110100001111110",
    "1110100110100101",
    "1110110100011000",
    "1111000111011000",
    "1111011011010100",
    "1111101101001001",
    "1111111011101111",
    "1111111000011110",
    "1111101110010110",
    "1111100100110100",
    "1111011011101101",
    "1111010011111100",
    "1111001111000100",
    "1111001110100110",
    "1111010011010111",
    "1111011100111000",
    "1111101001000101",
    "1111110101000001",
    "1111111101101010",
    "1111111111001100",
    "1111111101100111",
    "1111110101001000",
    "1111101001100101",
    "1111011101110011",
    "1111010100010011",
    "1111001110100011",
    "1111001101000010",
    "1111001111010111",
    "1111010100101111",
    "1111011100010100",
    "1111100101010011",
    "1111101111001000",
    "1111111001011101",
    "1111111011111011",
    "1111110001001110",
    "1111100110011011",
    "1111011011011110",
    "1111010000010100",
    "1111000101001101",
    "1110111011001010",
    "1110110011111011",
    "1110110001110001",
    "1110110110111001",
    "1111000100100101",
    "1111011010010100",
    "1111110101100000",
    "1111101110000101",
    "1111010101011010",
    "1111000100011101",
    "1110111101011001",
    "1110111111101100",
    "1111001000101101",
    "1111010100011101",
    "1111011111001000",
    "1111100110001011",
    "1111101001000100",
    "1111101001000101",
    "1111101000011111",
    "1111101001001011",
    "1111101011100101",
    "1111101110100011",
    "1111101111110000",
    "1111101101000000",
    "1111100101100000",
    "1111011010100010",
    "1111001111010111",
    "1111001000100010",
    "1111001010001110",
    "1111010110100100",
    "1111101100011011",
    "1111111000010001",
    "1111011101010110",
    "1111001000010001",
    "1110111100100001",
    "1110111010011110",
    "1110111111011110",
    "1111000111001011",
    "1111001101010100",
    "1111001111011001",
    "1111001101010111",
    "1111001001010101",
    "1111000110010110",
    "1111000111001001",
    "1111001100110111",
    "1111010110101000",
    "1111100001111101",
    "1111101011011111",
    "1111110000100100",
    "1111101111110110",
    "1111101001111101",
    "1111100000111000",
    "1111010111011000",
    "1111010000000101",
    "1111001100110010",
    "1111001110000010",
    "1111010011000011",
    "1111011010001001",
    "1111100001010101",
    "1111100111000010",
    "1111101010011101",
    "1111101011110011",
    "1111101011111111",
    "1111101100000110",
    "1111101100110011",
    "1111101101111101",
    "1111101110100100",
    "1111101101010111",
    "1111101001010101",
    "1111100010100100",
    "1111011010001111",
    "1111010010101100",
    "1111001110101001",
    "1111010000011100",
    "1111011001010110",
    "1111101001000000",
    "1111111101011010",
    "1111101100011111",
    "1111011000000100",
    "1111001000001001",
    "1110111110010100",
    "1110111010110111",
    "1110111100101010",
    "1111000001100111",
    "1111000111100111",
    "1111001100111000",
    "1111010000100100",
    "1111010010110001",
    "1111010100001011",
    "1111010101110001",
    "1111011000010001",
    "1111011011110011",
    "1111011111011110",
    "1111100001101011",
    "1111100000101100",
    "1111011011011011",
    "1111010010000000",
    "1111000110000001",
    "1110111010010001",
    "1110110001111110",
    "1110101111111111",
    "1110110101100111",
    "1111000010001010",
    "1111010011000101",
    "1111100100110100",
    "1111110100000011",
    "1111111110100100",
    "1111111100000101",
    "1111111010111111",
    "1111111100010000",
    "1111111110001100",
    "1111111111111100",
    "1111111110001110",
    "1111111011011010",
    "1111110110011000",
    "1111101110010010",
    "1111100010111110",
    "1111010101010000",
    "1111000110101000",
    "1110111001000110",
    "1110101110100011",
    "1110101000011101",
    "1110100111010101",
    "1110101010101111",
    "1110110001010111",
    "1110111001010101",
    "1111000000101100",
    "1111000110001110",
    "1111001001011101",
    "1111001010111101",
    "1111001011111100",
    "1111001101101101",
    "1111010001010010",
    "1111010110111011",
    "1111011110000101",
    "1111100101100010",
    "1111101011110001",
    "1111101111011100",
    "1111101111110001",
    "1111101100101000",
    "1111100110101100",
    "1111011111000111",
    "1111010111010101",
    "1111010000101100",
    "1111001100010100",
    "1111001010111111",
    "1111001101000100",
    "1111010010010101",
    "1111011010000100",
    "1111100011000000",
    "1111101011101110",
    "1111110011001001",
    "1111111000101111",
    "1111111100100110",
    "1111111111000101",
    "1111111111011001",
    "1111111110111010",
    "1111111111111011",
    "1111111100001001",
    "1111110100101001",
    "1111101001000010",
    "1111011010001100",
    "1111001010001110",
    "1110111100000111",
    "1110110010111011",
    "1110110001000010",
    "1110110111001101",
    "1111000100010111",
    "1111010101100101",
    "1111100111010101",
    "1111110110010011",
    "1111111111010011",
    "1111111001101011",
    "1111110111010010",
    "1111110101110000",
    "1111110010110111",
    "1111101101100010",
    "1111100110001110",
    "1111011110110001",
    "1111011001011110",
    "1111011000011010",
    "1111011100011100",
    "1111100101010011",
    "1111110001011000",
    "1111111110010111",
    "1111110110000010",
    "1111101101101011",
    "1111101001001010",
    "1111101000000010",
    "1111101001000110",
    "1111101011000001",
    "1111101100111110",
    "1111101111000001",
    "1111110010000100",
    "1111110111011011",
    "1111111111111000",
    "1111110011111101",
    "1111100110001000",
    "1111011000101101",
    "1111001110001111",
    "1111001000101010",
    "1111001000101000",
    "1111001101011110",
    "1111010101011011",
    "1111011110011110",
    "1111100110111110",
    "1111101110001011",
    "1111110100001010",
    "1111111001100101",
    "1111111111001000",
    "1111111010111101",
    "1111110101001011",
    "1111110000100000",
    "1111101110000001",
    "1111101110101001",
    "1111110010101111",
    "1111111010000110",
    "1111111100001010",
    "1111110001100010",
    "1111100111110101",
    "1111100000111000",
    "1111011110001010",
    "1111100000011010",
    "1111100111011011",
    "1111110010000111",
    "1111111110101100",
    "1111110100101101",
    "1111101001110000",
    "1111100001010010",
    "1111011011100110",
    "1111011000011011",
    "1111010111100000",
    "1111011000101000",
    "1111011100000001",
    "1111100010000011",
    "1111101011000101",
    "1111110110110010",
    "1111111100000010",
    "1111101111101001",
    "1111100110100101",
    "1111100011000011",
    "1111100110001000",
    "1111101111011000",
    "1111111100101111",
    "1111110100110111",
    "1111101000101010",
    "1111100000110001",
    "1111011101110000",
    "1111011110011111",
    "1111100000110110",
    "1111100010101100",
    "1111100010110100",
    "1111100001011010",
    "1111011111110110",
    "1111100000000011",
    "1111100011100010",
    "1111101010100001",
    "1111110011011100",
    "1111111011011110",
    "1111111111100001",
    "1111111101100000",
    "1111110101010001",
    "1111101000101111",
    "1111011011011000",
    "1111010001001010",
    "1111001101001111",
    "1111010001001101",
    "1111011100100101",
    "1111101101010100",
    "1111111111011111",
    "1111101100110100",
    "1111011100110101",
    "1111010000011100",
    "1111000111010101",
    "1111000000010010",
    "1110111010001001",
    "1110110100011101",
    "1110101111110011",
    "1110101101101110",
    "1110101111111101",
    "1110110111101000",
    "1111000100011100",
    "1111010100010010",
    "1111100011110001",
    "1111101111001100",
    "1111110011111101",
    "1111110001110100",
    "1111101011001001",
    "1111100100000110",
    "1111100000111101",
    "1111100100001101",
    "1111101101101000",
    "1111111010010011",
    "1111111010000101",
    "1111110011100100",
    "1111110100000000",
    "1111111010010111",
    "1111111100110001",
    "1111110101110111",
    "1111110100010111",
    "1111111001100101",
    "1111111011101000",
    "1111101110010101",
    "1111100010000011",
    "1111011001101011",
    "1111010110100100",
    "1111011000100000",
    "1111011110010110",
    "1111100110011111",
    "1111101111110010",
    "1111111001101010",
    "1111111011101000",
    "1111101111011110",
    "1111100001000101",
    "1111010000011111",
    "1110111111000010",
    "1110101111010110",
    "1110100100011111",
    "1110100001001100",
    "1110100110100000",
    "1110110011100001",
    "1111000101001000",
    "1111010111001001",
    "1111100101011011",
    "1111101101001001",
    "1111101101100110",
    "1111101000010000",
    "1111011111110110",
    "1111010111010001",
    "1111010000010010",
    "1111001011000111",
    "1111000110101010",
    "1111000001010010",
    "1110111001110000",
    "1110110000000000",
    "1110100101001101",
    "1110011011001111",
    "1110010100010010",
    "1110010010000011",
    "1110010101100100",
    "1110011110111011",
    "1110101101100001",
    "1111000000000111",
    "1111010101000110",
    "1111101010100111",
    "1111111110101011",
    "1111110000100110",
    "1111100100110111",
    "1111011110111010",
    "1111011110101000",
    "1111100010111101",
    "1111101010010000",
    "1111110010110000",
    "1111111010111111",
    "1111111101111000",
    "1111111000001101",
    "1111110100000111",
    "1111110001111011",
    "1111110010010001",
    "1111110101110110",
    "1111111100111100",
    "1111111000110000",
    "1111101100011011",
    "1111011111110011",
    "1111010101000000",
    "1111001101111011",
    "1111001011111100",
    "1111001111010001",
    "1111010111010000",
    "1111100010011100",
    "1111101111001000",
    "1111111011101111",
    "1111111000110010",
    "1111101110110011",
    "1111100101111011",
    "1111011101011011",
    "1111010100101100",
    "1111001011110000",
    "1111000011011010",
    "1110111101000010",
    "1110111010000001",
    "1110111011000100",
    "1110111111111011",
    "1111000111000011",
    "1111001110000100",
    "1111010010100100",
    "1111010010110100",
    "1111001110100110",
    "1111000111001001",
    "1110111110110001",
    "1110111000010000",
    "1110110101101010",
    "1110111000000100",
    "1110111111000000",
    "1111001000110100",
    "1111010011010111",
    "1111011100100011",
    "1111100011001111",
    "1111100111011100",
    "1111101010011000",
    "1111101101111001",
    "1111110011111010",
    "1111111101100011",
    "1111110101011000",
    "1111100110100100",
    "1111011000100011",
    "1111001110000000",
    "1111001000100111",
    "1111001000011101",
    "1111001011111101",
    "1111010000101110",
    "1111010100011100",
    "1111010110000000",
    "1111010110001000",
    "1111010111000011",
    "1111011011100110",
    "1111100101110010",
    "1111110101101101",
    "1111110110110111",
    "1111100011101111",
    "1111010101000000",
    "1111001101100100",
    "1111001110011100",
    "1111010110011000",
    "1111100010110001",
    "1111110000110001",
    "1111111110010000",
    "1111110101100111",
    "1111101010101011",
    "1111100000000101",
    "1111010101001101",
    "1111001010000100",
    "1110111111100001",
    "1110110110111111",
    "1110110010001000",
    "1110110010000101",
    "1110110111010001",
    "1111000001001000",
    "1111001110000111",
    "1111011011111000",
    "1111100111101001",
    "1111101110110111",
    "1111110000001000",
    "1111101011101001",
    "1111100011010101",
    "1111011010010001",
    "1111010011110001",
    "1111010010011001",
    "1111010111001011",
    "1111100001010100",
    "1111101110100101",
    "1111111100001010",
    "1111111000010011",
    "1111110000001010",
    "1111101011010010",
    "1111101000100110",
    "1111100110101010",
    "1111100100010101",
    "1111100001001100",
    "1111011101100100",
    "1111011010010011",
    "1111011000010001",
    "1111011000001000",
    "1111011010000111",
    "1111011110001100",
    "1111100100001010",
    "1111101011100101",
    "1111110100000000",
    "1111111100111010",
    "1111111010000110",
    "1111110001010010",
    "1111101000100011",
    "1111011111100100",
    "1111010110000000",
    "1111001011111111",
    "1111000010010000",
    "1110111010010011",
    "1110110101110001",
    "1110110101110111",
    "1110111010101111",
    "1111000011000011",
    "1111001100010100",
    "1111010011110100",
    "1111010111101100",
    "1111010111110010",
    "1111010110000011",
    "1111010101011101",
    "1111011001000111",
    "1111100010101001",
    "1111110001011011",
    "1111111101001000",
    "1111101100110111",
    "1111100001001111",
    "1111011100001111",
    "1111011101110101",
    "1111100100000011",
    "1111101100000001",
    "1111110010111001",
    "1111110110111110",
    "1111111000000100",
    "1111110111010101",
    "1111110110110110",
    "1111111000101001",
    "1111111101110111",
    "1111111001101010",
    "1111101111101001",
    "1111100110011111",
    "1111100000100001",
    "1111011111000010",
    "1111100001100111",
    "1111100110010000",
    "1111101001110101",
    "1111101001011011",
    "1111100011011101",
    "1111011000101111",
    "1111001100000010",
    "1111000001011001",
    "1110111100011011",
    "1110111110111011",
    "1111001000001000",
    "1111010100110011",
    "1111100000101100",
    "1111101000011010",
    "1111101010100001",
    "1111101000010100",
    "1111100101001000",
    "1111100100111100",
    "1111101010100100",
    "1111110110010110",
    "1111111010000011",
    "1111101010110100",
    "1111100000001010",
    "1111011100111010",
    "1111100001011110",
    "1111101011111011",
    "1111111001000000",
    "1111111010100111",
    "1111110001000100",
    "1111101010011011",
    "1111100100110100",
    "1111011101011110",
    "1111010010010000",
    "1111000010101100",
    "1110110000011110",
    "1110011110110110",
    "1110010001110000",
    "1110001100100011",
    "1110010001000101",
    "1110011111000000",
    "1110110011110100",
    "1111001011100101",
    "1111100001111110",
    "1111110011100110",
    "1111111110100011",
    "1111111101000110",
    "1111111101101000",
    "1111111111100000",
    "1111111100101100",
    "1111111011000100",
    "1111111010010110",
    "1111111001001010",
    "1111110110000001",
    "1111110000011000",
    "1111101001001001",
    "1111100010101001",
    "1111011111110001",
    "1111100010101110",
    "1111101011111011",
    "1111111001011101",
    "1111111000100110",
    "1111101110111100",
    "1111101101001001",
    "1111110100011010",
    "1111111100101110",
    "1111101001111011",
    "1111010111011010",
    "1111001000110100",
    "1111000000000011",
    "1110111100110010",
    "1110111101000010",
    "1110111110010001",
    "1110111110011001",
    "1110111100100011",
    "1110111001001110",
    "1110110101110001",
    "1110110011111011",
    "1110110101001101",
    "1110111010100000",
    "1111000011110100",
    "1111010000001010",
    "1111011101110011",
    "1111101010110100",
    "1111110101100111",
    "1111111101101000",
    "1111111100011110",
    "1111110110111110",
    "1111101111011100",
    "1111100100000000",
    "1111010100010000",
    "1111000001100001",
    "1110101110100001",
    "1110011110010100",
    "1110010011001101",
    "1110001110000111",
    "1110001110010010",
    "1110010010000000",
    "1110010111010101",
    "1110011101001001",
    "1110100011011101",
    "1110101011100110",
    "1110110111100010",
    "1111001001000110",
    "1111100000110000",
    "1111111100111000",
    "1111100101111110",
    "1111001100010011",
    "1110111010000001",
    "1110110001100001",
    "1110110010111110",
    "1110111100101011",
    "1111001011110011",
    "1111011101010111",
    "1111101110111011",
    "1111111110101101",
    "1111110100001111",
    "1111101010100100",
    "1111100100010101",
    "1111100001010010",
    "1111100001000011",
    "1111100011001111",
    "1111100111110010",
    "1111101110110100",
    "1111111000011011",
    "1111111011110001",
    "1111101111000010",
    "1111100011001011",
    "1111011010100000",
    "1111010111001011",
    "1111011010100110",
    "1111100100110011",
    "1111110100010010",
    "1111111001101010",
    "1111101000100001",
    "1111011011010011",
    "1111010011111110",
    "1111010011000101",
    "1111010111100111",
    "1111011111011111",
    "1111101000011100",
    "1111110000100111",
    "1111110111001110",
    "1111111100100000",
    "1111111110110000",
    "1111111001111110",
    "1111110101001011",
    "1111110001010110",
    "1111110000010000",
    "1111110011110111",
    "1111111101110000",
    "1111110001101101",
    "1111011011111111",
    "1111000100000000",
    "1110101101100011",
    "1110011100001111",
    "1110010010010010",
    "1110001111111011",
    "1110010011010101",
    "1110011001011000",
    "1110011110111010",
    "1110100001111101",
    "1110100010010010",
    "1110100001011010",
    "1110100010000010",
    "1110100110110010",
    "1110110001010000",
    "1111000001000101",
    "1111010011110011",
    "1111100101110100",
    "1111110011100101",
    "1111111010110011",
    "1111111010111111",
    "1111110101100100",
    "1111101101010001",
    "1111100101001000",
    "1111011111100001",
    "1111011101011100",
    "1111011110100110",
    "1111100001101110",
    "1111100101100000",
    "1111101001001101",
    "1111101100111110",
    "1111110001111000",
    "1111111001010111",
    "1111111011100001",
    "1111101101001011",
    "1111011101011100",
    "1111001111011010",
    "1111000110010010",
    "1111000100011000",
    "1111001010100011",
    "1111010111101010",
    "1111101001001100",
    "1111111011110101",
    "1111110011101110",
    "1111101000000010",
    "1111100010001101",
    "1111100001111101",
    "1111100101101110",
    "1111101011010111",
    "1111110000101111",
    "1111110100001010",
    "1111110100110001",
    "1111110010100011",
    "1111101110001000",
    "1111101000011111",
    "1111100010100110",
    "1111011100111111",
    "1111010111101101",
    "1111010010010111",
    "1111001100011100",
    "1111000101101110",
    "1110111110011011",
    "1110110111010001",
    "1110110001100001",
    "1110101110011001",
    "1110101111000010",
    "1110110011110110",
    "1110111100010111",
    "1111000111001000",
    "1111010001101100",
    "1111011001010110",
    "1111011011111010",
    "1111011000010110",
    "1111001111010111",
    "1111000011001010",
    "1110110110100111",
    "1110101100010110",
    "1110100101111001",
    "1110100011010111",
    "1110100011111011",
    "1110100110001110",
    "1110101001001100",
    "1110101100100110",
    "1110110001000000",
    "1110110111110100",
    "1111000010011111",
    "1111010001110110",
    "1111100101010111",
    "1111111010101110",
    "1111110001011000",
    "1111100010101111",
    "1111011011111101",
    "1111011101101001",
    "1111100110000011",
    "1111110001010000",
    "1111111010110101",
    "1111111111001100",
    "1111111100111111",
    "1111110101100001",
    "1111101011111010",
    "1111100011101111",
    "1111011111100100",
    "1111011111110110",
    "1111100010111011",
    "1111100101101111",
    "1111100101010000",
    "1111011111110000",
    "1111010101110111",
    "1111001010011000",
    "1111000001010000",
    "1110111110010111",
    "1111000011101001",
    "1111010000100110",
    "1111100010010111",
    "1111110100110100",
    "1111111011111001",
    "1111110010010011",
    "1111101110110011",
    "1111101111111001",
    "1111110011000111",
    "1111110101111111",
    "1111110111000001",
    "1111110101111010",
    "1111110011011101",
    "1111110000111100",
    "1111101111101000",
    "1111110000001101",
    "1111110010100101",
    "1111110110000010",
    "1111111001011101",
    "1111111011110011",
    "1111111100011100",
    "1111111011001101",
    "1111111000100011",
    "1111110101010011",
    "1111110010011101",
    "1111110001000000",
    "1111110001100101",
    "1111110100011001",
    "1111111001001001",
    "1111111111000011",
    "1111111010110111",
    "1111110101101011",
    "1111110001111100",
    "1111101111101011",
    "1111101110000111",
    "1111101011111110",
    "1111100111110000",
    "1111100000010101",
    "1111010101101010",
    "1111001000110000",
    "1110111011101011",
    "1110110000101110",
    "1110101001101111",
    "1110100111100010",
    "1110101001101010",
    "1110101110101011",
    "1110110100101111",
    "1110111010010011",
    "1110111110101011",
    "1111000010000010",
    "1111000101001011",
    "1111001000110010",
    "1111001100111100",
    "1111010000101001",
    "1111010010001111",
    "1111001111101011",
    "1111000111101101",
    "1110111010100101",
    "1110101010010100",
    "1110011010010001",
    "1110001110001101",
    "1110001001001110",
    "1110001100101101",
    "1110010111111001",
    "1110100111111111",
    "1110111001001001",
    "1111000111101101",
    "1111010001011001",
    "1111010110000011",
    "1111010111100101",
    "1111011000111110",
    "1111011100111100",
    "1111100100101001",
    "1111101111010000",
    "1111111010000101",
    "1111111110010011",
    "1111111100111101",
    "1111111100110100",
    "1111110000001001",
    "1111100000001100",
    "1111010001001100",
    "1111000111000110",
    "1111000100010010",
    "1111001000101111",
    "1111010010001010",
    "1111011100111101",
    "1111100101110110",
    "1111101011000111",
    "1111101101001101",
    "1111101110011111",
    "1111110001111001",
    "1111111001011110",
    "1111111010101000",
    "1111101100100000",
    "1111011111110001",
    "1111011000011011",
    "1111011001100011",
    "1111100100001010",
    "1111110110100001",
    "1111110011000101",
    "1111011101011100",
    "1111001100101010",
    "1111000011001111",
    "1111000001011111",
    "1111000101101100",
    "1111001100110111",
    "1111010011111000",
    "1111011000101101",
    "1111011010111101",
    "1111011011110000",
    "1111011100111111",
    "1111100000100011",
    "1111100111011000",
    "1111110001000010",
    "1111111011110000",
    "1111111011000011",
    "1111110110000000",
    "1111110110100100",
    "1111111100101001",
    "1111111001011100",
    "1111101110100001",
    "1111100101100101",
    "1111100000111110",
    "1111100001110110",
    "1111100111101110",
    "1111110000110000",
    "1111111010011000",
    "1111111101110000",
    "1111111001000110",
    "1111110111100111",
    "1111111000001001",
    "1111111001000010",
    "1111111000111000",
    "1111110111000101",
    "1111110100001101",
    "1111110001101111",
    "1111110001101000",
    "1111110101100000",
    "1111111101111101",
    "1111110101110001",
    "1111101000000010",
    "1111011011110101",
    "1111010100001010",
    "1111010011001011",
    "1111011001100111",
    "1111100110011110",
    "1111110111011000",
    "1111110110110011",
    "1111100111010010",
    "1111011100010011",
    "1111010110110010",
    "1111010110011011",
    "1111011001111101",
    "1111011111101110",
    "1111100110010010",
    "1111101101000000",
    "1111110011111100",
    "1111111011011111",
    "1111111100000111",
    "1111110011100010",
    "1111101100000100",
    "1111100111110001",
    "1111101000111010",
    "1111110001100011",
    "1111111101100010",
    "1111100101101111",
    "1111001010010110",
    "1110110000000011",
    "1110011011011101",
    "1110001111101110",
    "1110001101110010",
    "1110010100000110",
    "1110011111011111",
    "1110101100011011",
    "1110111000010000",
    "1111000001110001",
    "1111001001010000",
    "1111001111101000",
    "1111010101101100",
    "1111011011011011",
    "1111011111110110",
    "1111100001100001",
    "1111011111001101",
    "1111011000100010",
    "1111001110011001",
    "1111000010101100",
    "1110110111110100",
    "1110110000000101",
    "1110101101100001",
    "1110110001101110",
    "1110111101100110",
    "1111010000111011",
    "1111101010000101",
    "1111111001111110",
    "1111011111001100",
    "1111001001000110",
    "1110111010000111",
    "1110110010110011",
    "1110110001110011",
    "1110110100100100",
    "1110111000100000",
    "1110111011111010",
    "1110111110100100",
    "1111000001011110",
    "1111000101111001",
    "1111001100111000",
    "1111010110010000",
    "1111100000110000",
    "1111101010010000",
    "1111110000110000",
    "1111110011000101",
    "1111110001010011",
    "1111101100101100",
    "1111100111010010",
    "1111100011000011",
    "1111100001011010",
    "1111100010101110",
    "1111100110011001",
    "1111101011000100",
    "1111101111001011",
    "1111110001100001",
    "1111110001110011",
    "1111110000110100",
    "1111110000001001",
    "1111110001101100",
    "1111110111001000",
    "1111111110101011",
    "1111110000001001",
    "1111011110110110",
    "1111001101001111",
    "1110111110000000",
    "1110110011010111",
    "1110101110010001",
    "1110101110010100",
    "1110110001111110",
    "1110110111010110",
    "1110111100101110",
    "1111000001011010",
    "1111000101101001",
    "1111001010100101",
    "1111010001101100",
    "1111011100000010",
    "1111101001011100",
    "1111111000010110",
    "1111111001111011",
    "1111110000100001",
    "1111101101110010",
    "1111110010110011",
    "1111111110110110",
    "1111110000011001",
    "1111011110011110",
    "1111001111000100",
    "1111000101001101",
    "1111000010100001",
    "1111000110111110",
    "1111010001000000",
    "1111011110000111",
    "1111101011101100",
    "1111110111110111",
    "1111111101111101",
    "1111110101010101",
    "1111101100111111",
    "1111100011111001",
    "1111011001110100",
    "1111001111100001",
    "1111000110101010",
    "1111000001000111",
    "1111000000011001",
    "1111000101001101",
    "1111001110111000",
    "1111011011101011",
    "1111101001001011",
    "1111110101000000",
    "1111111101100111",
    "1111111101010011",
    "1111111010110101",
    "1111111001000010",
    "1111110101111010",
    "1111110000001000",
    "1111100111101110",
    "1111011110001111",
    "1111010110001001",
    "1111010010001000",
    "1111010011101111",
    "1111011010111100",
    "1111100101110001",
    "1111110001001010",
    "1111111001110101",
    "1111111101100111",
    "1111111011111101",
    "1111110110001011",
    "1111101110110000",
    "1111101000011000",
    "1111100100111100",
    "1111100100111011",
    "1111100111001110",
    "1111101001110111",
    "1111101010101101",
    "1111101000011011",
    "1111100011000110",
    "1111011100001111",
    "1111010110010000",
    "1111010011101001",
    "1111010110001110",
    "1111011110011110",
    "1111101011001011",
    "1111111001111101",
    "1111111000000110",
    "1111101101101101",
    "1111101000011110",
    "1111101000111001",
    "1111101110011010",
    "1111110111101110",
    "1111111100101010",
    "1111110000010010",
    "1111100100001110",
    "1111011001010110",
    "1111010000010001",
    "1111001001100010",
    "1111000101100101",
    "1111000100110100",
    "1111000111011101",
    "1111001101101101",
    "1111010111101100",
    "1111100101001000",
    "1111110101001010",
    "1111111001111111",
    "1111101010111100",
    "1111100000010100",
    "1111011100001010",
    "1111011111000111",
    "1111100111110101",
    "1111110011001101",
    "1111111101010011",
    "1111111101010011",
    "1111111110011110",
    "1111111010010111",
    "1111101111101111",
    "1111100101000101",
    "1111011101100110",
    "1111011011000111",
    "1111011101100110",
    "1111100011011010",
    "1111101001111100",
    "1111101110110001",
    "1111110000011011",
    "1111101110111001",
    "1111101011100001",
    "1111101000100100",
    "1111101000011000",
    "1111101100101010",
    "1111110101110110",
    "1111111101001011",
    "1111101110111001",
    "1111100010001000",
    "1111011001010110",
    "1111010101101010",
    "1111010110011011",
    "1111011001011101",
    "1111011011111101",
    "1111011011101010",
    "1111010111101101",
    "1111010001000010",
    "1111001001110100",
    "1111000100100111",
    "1111000011010111",
    "1111000110011011",
    "1111001100100110",
    "1111010011100010",
    "1111011000110100",
    "1111011010110101",
    "1111011001100011",
    "1111010110010101",
    "1111010011100001",
    "1111010011111011",
    "1111011001111101",
    "1111100110110110",
    "1111111001110110",
    "1111101111101011",
    "1111011001101011",
    "1111001000000100",
    "1110111101101101",
    "1110111011101010",
    "1111000001000011",
    "1111001011100101",
    "1111011000011101",
    "1111100101011011",
    "1111110001011100",
    "1111111100011010",
    "1111111001001011",
    "1111101111000101",
    "1111100101011111",
    "1111011101001110",
    "1111010111010110",
    "1111010100110111",
    "1111010110001000",
    "1111011010110100",
    "1111100001111101",
    "1111101010010101",
    "1111110010110110",
    "1111111010100011",
    "1111111111001110",
    "1111111011000110",
    "1111111001001000",
    "1111111000111100",
    "1111111001110000",
    "1111111010100001",
    "1111111010010100",
    "1111111000101000",
    "1111110101100110",
    "1111110001111100",
    "1111101110110011",
    "1111101101010101",
    "1111101110001000",
    "1111110000111010",
    "1111110100100100",
    "1111110111011011",
    "1111110111111000",
    "1111110100111110",
    "1111101110111111",
    "1111100111011000",
    "1111100000010111",
    "1111011100001100",
    "1111011100010100",
    "1111100000111110",
    "1111101001000110",
    "1111110010100111",
    "1111111011000101",
    "1111111111100101",
    "1111111110101000",
    "1111111110010000",
    "1111111000101110",
    "1111110011001010",
    "1111101111111101",
    "1111110000100110",
    "1111110101001000",
    "1111111011111010",
    "1111111101110110",
    "1111111011011001",
    "1111111111000011",
    "1111110110011000",
    "1111100110011000",
    "1111010100000101",
    "1111000011101001",
    "1110111000111111",
    "1110110110101111",
    "1110111101001111",
    "1111001010101101",
    "1111011011100101",
    "1111101011110010",
    "1111110111110110",
    "1111111101101111",
    "1111111101001011",
    "1111110111101100",
    "1111101111101011",
    "1111100111100001",
    "1111100000111001",
    "1111011100011110",
    "1111011010000010",
    "1111011000111110",
    "1111011000100111",
    "1111011000100011",
    "1111011000111001",
    "1111011010000111",
    "1111011100111100",
    "1111100001111001",
    "1111101001001011",
    "1111110010001001",
    "1111111011101111",
    "1111111011100010",
    "1111110101010001",
    "1111110010101000",
    "1111110100010001",
    "1111111010001110",
    "1111111100000100",
    "1111101111110011",
    "1111100010010101",
    "1111010101001011",
    "1111001001100011",
    "1111000000011001",
    "1110111001111100",
    "1110110101111110",
    "1110110011110100",
    "1110110010100100",
    "1110110001011110",
    "1110110000000111",
    "1110101110101000",
    "1110101101100001",
    "1110101101100011",
    "1110101111001100",
    "1110110010100111",
    "1110110111101000",
    "1110111101110000",
    "1111000100100000",
    "1111001011100101",
    "1111010010110110",
    "1111011010100000",
    "1111100011000000",
    "1111101100111011",
    "1111111000100010",
    "1111111010011010",
    "1111101100111110",
    "1111100000101011",
    "1111010111001000",
    "1111010001101100",
    "1111010000111101",
    "1111010100101110",
    "1111011100001001",
    "1111100110000011",
    "1111110000111000",
    "1111111011000011",
    "1111111100110110",
    "1111110111111100",
    "1111110110011101",
    "1111110111111100",
    "1111111011010010",
    "1111111111000110",
    "1111111110000001",
    "1111111101010111",
    "1111111111110000",
    "1111111010011010",
    "1111110001100101",
    "1111100110100101",
    "1111011010101000",
    "1111001110111010",
    "1111000100011010",
    "1110111011101011",
    "1110110101000000",
    "1110110000011001",
    "1110101101111010",
    "1110101101110010",
    "1110110000100011",
    "1110110110111111",
    "1111000001111000",
    "1111010001011001",
    "1111100100110001",
    "1111111010000011",
    "1111110001100011",
    "1111100001000010",
    "1111010110011010",
    "1111010010100001",
    "1111010100100101",
    "1111011011000001",
    "1111100011111100",
    "1111101110000111",
    "1111111001001000",
    "1111111010111001",
    "1111101101111110",
    "1111100000100100",
    "1111010011111011",
    "1111001001101010",
    "1111000011100010",
    "1111000010101001",
    "1111000111001001",
    "1111010000010001",
    "1111011100101000",
    "1111101010100101",
    "1111111000011000",
    "1111111011101011",
    "1111110011000011",
    "1111101110100100",
    "1111101110010010",
    "1111110001010111",
    "1111110110010001",
    "1111111011000010",
    "1111111101111011",
    "1111111101111100",
    "1111111010111111",
    "1111110101110011",
    "1111101111100100",
    "1111101001100011",
    "1111100100101001",
    "1111100001001111",
    "1111011111001101",
    "1111011110000000",
    "1111011100111000",
    "1111011011000100",
    "1111011000001000",
    "1111010011111000",
    "1111001110101000",
    "1111001001000111",
    "1111000100010000",
    "1111000000111110",
    "1111000000000111",
    "1111000010001010",
    "1111000111011000",
    "1111001111110001",
    "1111011010111100",
    "1111101000000111",
    "1111110110001001",
    "1111111100011000",
    "1111110001000101",
    "1111101001001011",
    "1111100101011011",
    "1111100110000011",
    "1111101010101000",
    "1111110010011011",
    "1111111100100001",
    "1111111000001000",
    "1111101100101001",
    "1111100010000101",
    "1111011001100010",
    "1111010011110110",
    "1111010001100001",
    "1111010010011010",
    "1111010101110100",
    "1111011010100000",
    "1111011111000100",
    "1111100010010000",
    "1111100011001010",
    "1111100001011001",
    "1111011100111010",
    "1111010101111001",
    "1111001100101010",
    "1111000001110001",
    "1110110110001101",
    "1110101011001001",
    "1110100001111110",
    "1110011011110101",
    "1110011001011110",
    "1110011011000100",
    "1110011111111101",
    "1110100111000110",
    "1110101111010001",
    "1110110111010101",
    "1110111110011100",
    "1111000100000000",
    "1111000111011010",
    "1111001000001001",
    "1111000101111011",
    "1111000000100110",
    "1110111000100111",
    "1110101110110110",
    "1110100100110110",
    "1110011100001010",
    "1110010110001110",
    "1110010011111001",
    "1110010101010111",
    "1110011010010001",
    "1110100001110110",
    "1110101011001010",
    "1110110101010010",
    "1110111111011110",
    "1111001001010000",
    "1111010010001101",
    "1111011010000010",
    "1111100000100011",
    "1111100101100101",
    "1111101001010000",
    "1111101011110111",
    "1111101101111010",
    "1111110000000001",
    "1111110010101101",
    "1111110110010000",
    "1111111010101011",
    "1111111111111000",
    "1111111010010010",
    "1111110100000010",
    "1111101101011011",
    "1111100110110011",
    "1111100000100110",
    "1111011011100011",
    "1111011000010110",
    "1111010111100000",
    "1111011001000010",
    "1111011100101000",
    "1111100001111001",
    "1111101000101110",
    "1111110001001010",
    "1111111011001101",
    "1111111001110101",
    "1111101111110001",
    "1111101001001000",
    "1111101000100101",
    "1111101111011111",
    "1111111100111001",
    "1111110010101010",
    "1111100100010011",
    "1111011101000100",
    "1111100000000010",
    "1111101101001000",
    "1111111111000011",
    "1111101001111111",
    "1111011000111001",
    "1111001110111000",
    "1111001100010011",
    "1111001110111111",
    "1111010011101111",
    "1111011000000011",
    "1111011010110010",
    "1111011100010111",
    "1111011101110111",
    "1111011111111010",
    "1111100010010111",
    "1111100100011010",
    "1111100101000110",
    "1111100100000011",
    "1111100001111101",
    "1111100000001101",
    "1111100000011111",
    "1111100011111001",
    "1111101010100011",
    "1111110011100001",
    "1111111101010111",
    "1111111001001011",
    "1111110000011010",
    "1111100111100011",
    "1111011101100001",
    "1111010001101100",
    "1111000100101100",
    "1110111000010000",
    "1110101110101110",
    "1110101010011000",
    "1110101100101010",
    "1110110101101010",
    "1111000100001000",
    "1111010101111110",
    "1111101000101011",
    "1111111001111101",
    "1111110111111000",
    "1111101110000000",
    "1111101000110010",
    "1111101000001100",
    "1111101100000001",
    "1111110100000000",
    "1111111111101010",
    "1111110010000011",
    "1111100011001010",
    "1111010110010010",
    "1111001110001010",
    "1111001100101010",
    "1111010010001011",
    "1111011101100110",
    "1111101100010101",
    "1111111011010100",
    "1111111000000110",
    "1111101111100100",
    "1111101011010010",
    "1111101010100001",
    "1111101100010101",
    "1111110000011001",
    "1111110111001110",
    "1111111110001110",
    "1111101111100101",
    "1111011101100110",
    "1111001010011110",
    "1110111001011000",
    "1110101101100000",
    "1110101001010101",
    "1110101101111010",
    "1110111010100011",
    "1111001100111010",
    "1111100001101100",
    "1111110101010111",
    "1111111010111000",
    "1111110000101110",
    "1111101100001110",
    "1111101100010110",
    "1111101111100001",
    "1111110100101001",
    "1111111011101100",
    "1111111010001110",
    "1111101011110010",
    "1111011000101000",
    "1111000010000101",
    "1110101011010011",
    "1110011000011110",
    "1110001101110000",
    "1110001101111000",
    "1110011001001100",
    "1110101101010100",
    "1111000101111001",
    "1111011101111011",
    "1111110001001111",
    "1111111101010100",
    "1111111110011010",
    "1111111110101101",
    "1111110110001010",
    "1111101001010011",
    "1111011001011000",
    "1111000111101101",
    "1110110101110110",
    "1110100101101100",
    "1110011001011001",
    "1110010010111101",
    "1110010011110100",
    "1110011100101101",
    "1110101101000111",
    "1111000011011100",
    "1111011100111101",
    "1111110110010111",
    "1111110011011111",
    "1111100011000000",
    "1111011001001110",
    "1111010110001101",
    "1111011001011011",
    "1111100010011100",
    "1111110000110111",
    "1111111100000010",
    "1111100101110100",
    "1111001110110101",
    "1110111001111111",
    "1110101010001100",
    "1110100001101011",
    "1110100001011001",
    "1110101001000110",
    "1110110111011111",
    "1111001010100011",
    "1111011111111000",
    "1111110100110111",
    "1111111000110100",
    "1111101011001010",
    "1111100011100010",
    "1111100010101110",
    "1111101000101101",
    "1111110100101001",
    "1111111011000001",
    "1111101000011000",
    "1111010101100010",
    "1111000100100010",
    "1110110111001000",
    "1110101110101101",
    "1110101100011011",
    "1110110001001010",
    "1110111101010100",
    "1111010000100001",
    "1111101001001101",
    "1111111011011001",
    "1111100001000010",
    "1111001011010001",
    "1110111100110101",
    "1110110110110110",
    "1110111000101100",
    "1111000000100001",
    "1111001100001100",
    "1111011010000001",
    "1111101001001100",
    "1111111001100001",
    "1111110101001010",
    "1111100011110001",
    "1111010100000110",
    "1111001000100111",
    "1111000011111001",
    "1111000111110010",
    "1111010100110011",
    "1111101001101101",
    "1111111100001001",
    "1111100000010111",
    "1111000110011010",
    "1110110001000011",
    "1110100001111011",
    "1110011001100011",
    "1110010111100011",
    "1110011011001010",
    "1110100011110100",
    "1110110001010010",
    "1111000011011100",
    "1111011001111010",
    "1111110011001011",
    "1111110011100110",
    "1111011110010111",
    "1111010001000111",
    "1111001110101011",
    "1111010111101101",
    "1111101010100001",
    "1111111100101100",
    "1111100010100010",
    "1111001011001001",
    "1110111001010110",
    "1110101110100011",
    "1110101011001001",
    "1110101111001111",
    "1110111010110100",
    "1111001101100000",
    "1111100110000011",
    "1111111101111011",
    "1111100010001101",
    "1111001010110101",
    "1110111011011110",
    "1110110110011000",
    "1110111011111100",
    "1111001010110101",
    "1111100000101100",
    "1111111010101110",
    "1111101001110110",
    "1111001111101110",
    "1110111001001001",
    "1110100111111001",
    "1110011101001010",
    "1110011001100011",
    "1110011101000100",
    "1110100111010001",
    "1110110111101100",
    "1111001101010100",
    "1111100110011101",
    "1111111111100010",
    "1111101000010010",
    "1111010111101100",
    "1111010001010100",
    "1111010111000100",
    "1111101000011000",
    "1111111101111111",
    "1111100001001010",
    "1111000110100000",
    "1110110010001101",
    "1110100110011010",
    "1110100011000101",
    "1110100110110100",
    "1110110000000111",
    "1110111110010100",
    "1111010001101001",
    "1111101010001111",
    "1111111000111111",
    "1111011011000010",
    "1111000000001000",
    "1110101100110010",
    "1110100100010011",
    "1110100111110101",
    "1110110110001000",
    "1111001011111010",
    "1111100101001011",
    "1111111110001100",
    "1111101011101001",
    "1111011001110111",
    "1111001101000010",
    "1111000101100111",
    "1111000100001110",
    "1111001001111010",
    "1111010111011101",
    "1111101100011100",
    "1111111001001001",
    "1111011100111100",
    "1111000011000110",
    "1110101111010111",
    "1110100100000001",
    "1110100001011111",
    "1110100110011101",
    "1110110000100111",
    "1110111101010111",
    "1111001010011000",
    "1111010110000110",
    "1111011111101110",
    "1111100111000101",
    "1111101100001101",
    "1111101111000101",
    "1111101111100000",
    "1111101101010010",
    "1111101000011101",
    "1111100001011100",
    "1111011001010001",
    "1111010001011111",
    "1111001100000100",
    "1111001011010011",
    "1111010001011100",
    "1111100000000010",
    "1111110110111010",
    "1111101100010100",
    "1111001101110101",
    "1110110010001101",
    "1110011101001001",
    "1110010000010111",
    "1110001011101000",
    "1110001101001110",
    "1110010011001011",
    "1110011100100000",
    "1110101001001110",
    "1110111001111100",
    "1111001110110011",
    "1111100110101101",
    "1111111111000110",
    "1111101011010110",
    "1111011011111111",
    "1111010100110110",
    "1111010110010000",
    "1111011110111000",
    "1111101100011001",
    "1111111100001100",
    "1111110011111010",
    "1111100101011000",
    "1111011001000110",
    "1111001111101000",
    "1111001001011101",
    "1111000110111110",
    "1111001000011000",
    "1111001101110010",
    "1111010111000011",
    "1111100011100010",
    "1111110010001010",
    "1111111110100100",
    "1111110000011011",
    "1111100101000001",
    "1111011101101001",
    "1111011011000100",
    "1111011101010100",
    "1111100011100100",
    "1111101100001011",
    "1111110101001111",
    "1111111101000011",
    "1111111101010100",
    "1111111010001000",
    "1111111001000011",
    "1111111001110000",
    "1111111100010110",
    "1111111110101010",
    "1111110110110100",
    "1111101100001010",
    "1111011111101100",
    "1111010011011000",
    "1111001001100011",
    "1111000100001110",
    "1111000100100101",
    "1111001010100110",
    "1111010101000110",
    "1111100010010100",
    "1111110000011101",
    "1111111110010100",
    "1111110100101000",
    "1111101000100011",
    "1111011101011110",
    "1111010011111100",
    "1111001101000000",
    "1111001010000001",
    "1111001011110111",
    "1111010010100001",
    "1111011100100110",
    "1111100111011111",
    "1111110000000111",
    "1111110011111100",
    "1111110001101010",
    "1111101001100101",
    "1111011101010010",
    "1111001111001010",
    "1111000001011111",
    "1110110101111011",
    "1110101101010111",
    "1110101000001100",
    "1110100110100101",
    "1110101001000100",
    "1110110000100100",
    "1110111110010010",
    "1111010010110011",
    "1111101101001111",
    "1111110100110011",
    "1111010111001000",
    "1110111101110011",
    "1110101100010100",
    "1110100100011101",
    "1110100110000011",
    "1110101111010111",
    "1110111101101011",
    "1111001110001111",
    "1111011110101101",
    "1111101101001111",
    "1111111000101001",
    "1111111111101010",
    "1111111011111101",
    "1111111100000111",
    "1111111111110001",
    "1111111001100110",
    "1111110000111011",
    "1111100111010100",
    "1111011110001001",
    "1111010110110111",
    "1111010010111101",
    "1111010011011100",
    "1111011000110111",
    "1111100011000011",
    "1111110000110010",
    "1111111111110001",
    "1111110000111011",
    "1111100100100111",
    "1111011100000101",
    "1111010111110010",
    "1111010111010101",
    "1111011010001001",
    "1111011111100110",
    "1111100111011011",
    "1111110001011000",
    "1111111100111100",
    "1111110111000100",
    "1111101100101010",
    "1111100110010110",
    "1111100110100100",
    "1111101110101101",
    "1111111110011101",
    "1111101100011000",
    "1111010101011010",
    "1111000000011001",
    "1110110000010001",
    "1110100110011111",
    "1110100010111000",
    "1110100100001110",
    "1110101001001001",
    "1110110000100110",
    "1110111010000111",
    "1111000101100010",
    "1111010010011100",
    "1111011111110101",
    "1111101011111110",
    "1111110100110101",
    "1111111000101101",
    "1111110110111011",
    "1111110000001100",
    "1111100110100101",
    "1111011100111000",
    "1111010110000001",
    "1111010100010010",
    "1111011000111010",
    "1111100011101111",
    "1111110011011011",
    "1111111010001100",
    "1111100111101101",
    "1111010111010011",
    "1111001010100011",
    "1111000010001011",
    "1110111110011110",
    "1110111111100011",
    "1111000101011111",
    "1111001111111011",
    "1111011101100110",
    "1111101100011110",
    "1111111010000011",
    "1111111011101110",
    "1111110110000110",
    "1111110100110111",
    "1111110110101101",
    "1111111001111000",
    "1111111100111001",
    "1111111111001001",
    "1111111111000010",
    "1111111100111100",
    "1111111001110001",
    "1111110101001111",
    "1111101111110100",
    "1111101010101011",
    "1111100111001001",
    "1111100110011000",
    "1111101000110111",
    "1111101110010110",
    "1111110110000010",
    "1111111110110000",
    "1111111000101011",
    "1111110001011111",
    "1111101100100011",
    "1111101010011010",
    "1111101011001010",
    "1111101110100010",
    "1111110011111111",
    "1111111010110100",
    "1111111101101011",
    "1111110110001100",
    "1111101111010100",
    "1111101001100000",
    "1111100101001011",
    "1111100010100110",
    "1111100001111110",
    "1111100011010000",
    "1111100110000110",
    "1111101001110011",
    "1111101101011001",
    "1111101111110110",
    "1111110000011110",
    "1111101111001000",
    "1111101100011110",
    "1111101001101101",
    "1111101000001111",
    "1111101001000110",
    "1111101100100111",
    "1111110010010000",
    "1111111000110111",
    "1111111111000101",
    "1111111100010000",
    "1111111001111001",
    "1111111001111000",
    "1111111011110110",
    "1111111111001010",
    "1111111100100110",
    "1111110111110010",
    "1111110010010010",
    "1111101011111000",
    "1111100100010111",
    "1111011011110111",
    "1111010011000000",
    "1111001010101111",
    "1111000011111110",
    "1110111111011111",
    "1110111101101011",
    "1110111110011100",
    "1111000001100010",
    "1111000110101000",
    "1111001101011100",
    "1111010101101111",
    "1111011111000111",
    "1111101000111000",
    "1111110001110110",
    "1111111000100111",
    "1111111011101001",
    "1111111001110100",
    "1111110010110000",
    "1111100111001001",
    "1111011000101100",
    "1111001001110010",
    "1110111100110101",
    "1110110011110001",
    "1110101111100011",
    "1110101111110110",
    "1110110011100010",
    "1110111000110111",
    "1110111110000111",
    "1111000010001011",
    "1111000100110011",
    "1111000110011011",
    "1111001000000100",
    "1111001010101111",
    "1111001111001010",
    "1111010101100000",
    "1111011101010001",
    "1111100101011111",
    "1111101100111011",
    "1111110010011010",
    "1111110101001110",
    "1111110101001011",
    "1111110010110110",
    "1111101111011000",
    "1111101100010000",
    "1111101010111010",
    "1111101100010111",
    "1111110001000001",
    "1111111000100101",
    "1111111101101001",
    "1111110010110011",
    "1111100111111010",
    "1111011101111000",
    "1111010101001110",
    "1111001110010001",
    "1111001001001001",
    "1111000110000100",
    "1111000101011101",
    "1111000111110101",
    "1111001101111101",
    "1111011000011011",
    "1111100111001001",
    "1111111001001001",
    "1111110011100001",
    "1111100001100100",
    "1111010011100010",
    "1111001011100000",
    "1111001010011110",
    "1111010000011001",
    "1111011100100000",
    "1111101101011010",
    "1111111110101001",
    "1111101001111111",
    "1111010111010001",
    "1111001001010000",
    "1111000010001000",
    "1111000011001010",
    "1111001100001111",
    "1111011011111000",
    "1111101111110110",
    "1111111010011101",
    "1111100101100101",
    "1111010011011111",
    "1111000101011111",
    "1110111100010111",
    "1110111000011010",
    "1110111001011001",
    "1110111110110110",
    "1111000111111001",
    "1111010011011010",
    "1111100000011001",
    "1111101101110100",
    "1111111010110101",
    "1111111001010011",
    "1111101111011000",
    "1111101000000001",
    "1111100011110011",
    "1111100010111000",
    "1111100101000000",
    "1111101001010000",
    "1111101110011000",
    "1111110011001011",
    "1111110110111011",
    "1111111001100011",
    "1111111011011101",
    "1111111101010010",
    "1111111111100011",
    "1111111101101001",
    "1111111010110100",
    "1111111000101011",
    "1111111000001000",
    "1111111001110111",
    "1111111110001011",
    "1111111011000000",
    "1111110010000111",
    "1111100111011101",
    "1111011011001111",
    "1111001101101000",
    "1110111110111101",
    "1110110000001000",
    "1110100010011101",
    "1110010111010101",
    "1110001111111000",
    "1110001100011110",
    "1110001100101110",
    "1110001111101110",
    "1110010100100010",
    "1110011010100000",
    "1110100001100010",
    "1110101010000100",
    "1110110100101001",
    "1111000001110001",
    "1111010001011111",
    "1111100011000000",
    "1111110100101111",
    "1111111011010111",
    "1111101111100000",
    "1111101001000101",
    "1111101000100101",
    "1111101101010001",
    "1111110101011110",
    "1111111111001100",
    "1111110111011010",
    "1111101111101100",
    "1111101010001010",
    "1111100110110110",
    "1111100101101001",
    "1111100110100011",
    "1111101001111101",
    "1111110000010001",
    "1111111001100100",
    "1111111010100110",
    "1111101101100100",
    "1111100000111101",
    "1111010110100000",
    "1111001111011111",
    "1111001100011001",
    "1111001101000100",
    "1111010000111011",
    "1111010111001110",
    "1111011111010110",
    "1111101000111111",
    "1111110100000101",
    "1111111111010110",
    "1111110001101101",
    "1111100011110011",
    "1111010110110010",
    "1111001100000101",
    "1111000100110001",
    "1111000001001111",
    "1111000001001101",
    "1111000011101100",
    "1111000111011101",
    "1111001011001110",
    "1111001101111101",
    "1111001111000111",
    "1111001110101001",
    "1111001100101110",
    "1111001001110010",
    "1111000110001110",
    "1111000010010101",
    "1110111110010010",
    "1110111010001110",
    "1110110110010011",
    "1110110010101100",
    "1110101111101000",
    "1110101101010111",
    "1110101100001100",
    "1110101100010110",
    "1110101101111101",
    "1110110001000101",
    "1110110101100111",
    "1110111011011101",
    "1111000010100100",
    "1111001011000010",
    "1111010100111110",
    "1111100000010100",
    "1111101100100110",
    "1111111001000100",
    "1111111011010001",
    "1111110001011101",
    "1111101010010001",
    "1111100110001000",
    "1111100101000001",
    "1111100110101101",
    "1111101010101101",
    "1111110000011100",
    "1111110111001011",
    "1111111101111101",
    "1111111100001110",
    "1111111000101100",
    "1111111000011111",
    "1111111100010111",
    "1111111011100100",
    "1111110000000001",
    "1111100010011010",
    "1111010100101010",
    "1111001000110010",
    "1111000000011010",
    "1110111100101011",
    "1110111101110011",
    "1111000011010000",
    "1111001011110010",
    "1111010101101111",
    "1111011111101011",
    "1111101000100101",
    "1111110000001000",
    "1111110110101000",
    "1111111100101110",
    "1111111100111011",
    "1111110110001101",
    "1111101111010111",
    "1111101001000101",
    "1111100100010101",
    "1111100001111110",
    "1111100010011111",
    "1111100101111110",
    "1111101100000100",
    "1111110100000010",
    "1111111100111101",
    "1111111010000110",
    "1111110010000110",
    "1111101011111001",
    "1111101000001111",
    "1111100111100111",
    "1111101010000010",
    "1111101110111110",
    "1111110101100010",
    "1111111100101001",
    "1111111100100000",
    "1111110110011010",
    "1111110001000111",
    "1111101100011110",
    "1111101000010111",
    "1111100100110111",
    "1111100010011001",
    "1111100001010101",
    "1111100010001101",
    "1111100101010000",
    "1111101010011100",
    "1111110001100111",
    "1111111010011101",
    "1111111011001001",
    "1111101111011011",
    "1111100010100001",
    "1111010100110111",
    "1111000111011111",
    "1110111011101101",
    "1110110011001000",
    "1110101110111010",
    "1110101111101001",
    "1110110101000110",
    "1110111110001100",
    "1111001001011001",
    "1111010101001011",
    "1111011111111011",
    "1111101000100001",
    "1111101110000000",
    "1111101111111101",
    "1111101110010100",
    "1111101001010111",
    "1111100001110001",
    "1111011000011110",
    "1111001110101110",
    "1111000101101110",
    "1110111110011100",
    "1110111001100011",
    "1110110111000110",
    "1110110110110001",
    "1110110111111110",
    "1110111010001001",
    "1110111100111000",
    "1111000000000000",
    "1111000011101010",
    "1111001000001011",
    "1111001101110011",
    "1111010100100100",
    "1111011100000010",
    "1111100011010101",
    "1111101001010001",
    "1111101100101111",
    "1111101101000101",
    "1111101010011001",
    "1111100101100000",
    "1111011111111111",
    "1111011011100001",
    "1111011001111001",
    "1111011100010111",
    "1111100011011101",
    "1111101110101111",
    "1111111100101100",
    "1111110100101110",
    "1111100111111000",
    "1111011110101000",
    "1111011010000110",
    "1111011010100011",
    "1111011111100100",
    "1111101000001010",
    "1111110011001011",
    "1111111111001111",
    "1111110101000111",
    "1111101011010101",
    "1111100100100010",
    "1111100001010010",
    "1111100001100001",
    "1111100100010111",
    "1111101000010111",
    "1111101011111000",
    "1111101101011111",
    "1111101100100000",
    "1111101001000111",
    "1111100100011010",
    "1111100000000010",
    "1111011101110010",
    "1111011111000010",
    "1111100100100000",
    "1111101110000111",
    "1111111010110011",
    "1111110111001001",
    "1111101001111101",
    "1111011111110000",
    "1111011010000100",
    "1111011001100101",
    "1111011101111010",
    "1111100101110100",
    "1111101111100010",
    "1111111001011000",
    "1111111101110101",
    "1111110110111110",
    "1111110010010011",
    "1111110000000000",
    "1111110000001111",
    "1111110011001000",
    "1111111000101101",
    "1111111111011101",
    "1111110110011011",
    "1111101101101010",
    "1111100110110010",
    "1111100011001011",
    "1111100011100001",
    "1111100111101101",
    "1111101111001000",
    "1111111000101101",
    "1111111100110010",
    "1111110010101100",
    "1111101010001110",
    "1111100100100010",
    "1111100010011101",
    "1111100100011000",
    "1111101001111011",
    "1111110010000011",
    "1111111011001000",
    "1111111100100110",
    "1111110110101110",
    "1111110100000011",
    "1111110100100111",
    "1111110111100111",
    "1111111011110100",
    "1111111111111001",
    "1111111101001110",
    "1111111100010011",
    "1111111101101011",
    "1111111110010101",
    "1111110111101110",
    "1111101110101011",
    "1111100011111001",
    "1111011000100010",
    "1111001110000010",
    "1111000101110110",
    "1111000000111110",
    "1110111111110000",
    "1111000001110001",
    "1111000110010000",
    "1111001100010001",
    "1111010011000101",
    "1111011010010001",
    "1111100001100110",
    "1111101000111100",
    "1111110000001001",
    "1111110111000001",
    "1111111101011010",
    "1111111100100011",
    "1111110110101111",
    "1111110000110110",
    "1111101010111001",
    "1111100101010011",
    "1111100000111101",
    "1111011110111010",
    "1111100000001101",
    "1111100101011011",
    "1111101110011000",
    "1111111001111110",
    "1111111001101001",
    "1111101110111101",
    "1111101000011001",
    "1111100111111011",
    "1111101110101000",
    "1111111100010000",
    "1111110000111110",
    "1111011100000111",
    "1111001000101101",
    "1110111010000100",
    "1110110010011100",
    "1110110010110110",
    "1110111010110100",
    "1111001000111001",
    "1111011010110000",
    "1111101101101110",
    "1111111110111011",
    "1111110100011100",
    "1111101110110100",
    "1111110001011010",
    "1111111011110010",
    "1111110100010100",
    "1111100010100001",
    "1111010010101100",
    "1111000111110001",
    "1111000011001101",
    "1111000100110100",
    "1111001011010110",
    "1111010101011111",
    "1111100010011100",
    "1111110001111110",
    "1111111100000010",
    "1111101000100101",
    "1111010101011101",
    "1111000101000001",
    "1110111001011001",
    "1110110011110001",
    "1110110011111001",
    "1110111000011000",
    "1110111111001111",
    "1111000110100111",
    "1111001101001111",
    "1111010010011100",
    "1111010110000011",
    "1111011000001100",
    "1111011001001100",
    "1111011001100101",
    "1111011010000111",
    "1111011011110010",
    "1111011111100001",
    "1111100101101010",
    "1111101101110100",
    "1111110110100110",
    "1111111110001010",
    "1111111101001111",
    "1111111100110100",
    "1111111111001011",
    "1111110111100111",
    "1111101101111011",
    "1111100100000011",
    "1111011011111000",
    "1111010110111110",
    "1111010110010101",
    "1111011010010001",
    "1111100010011101",
    "1111101110000011",
    "1111111011110101",
    "1111110101011111",
    "1111100111011000",
    "1111011011000111",
    "1111010001111000",
    "1111001100100000",
    "1111001011010100",
    "1111001110001010",
    "1111010100010101",
    "1111011100110000",
    "1111100110001000",
    "1111101111001010",
    "1111110110101001",
    "1111111011110011",
    "1111111110010001",
    "1111111110001001",
    "1111111011111110",
    "1111111000100100",
    "1111110100110110",
    "1111110001110110",
    "1111110000100110",
    "1111110001111101",
    "1111110110010011",
    "1111111101010010",
    "1111111010001010",
    "1111110001110010",
    "1111101011010001",
    "1111100111111100",
    "1111101000010000",
    "1111101011101000",
    "1111110000101011",
    "1111110101100100",
    "1111111000101101",
    "1111111000110011",
    "1111110101001110",
    "1111101101110101",
    "1111100011001000",
    "1111010110001101",
    "1111001000100011",
    "1110111011111000",
    "1110110001110110",
    "1110101011100110",
    "1110101001100011",
    "1110101011010110",
    "1110110000000101",
    "1110110110110010",
    "1110111110101000",
    "1111000111010000",
    "1111010000100011",
    "1111011010011011",
    "1111100100100111",
    "1111101110011110",
    "1111110111001111",
    "1111111110000110",
    "1111111101001111",
    "1111111010100010",
    "1111111000110010",
    "1111110110110010",
    "1111110011100001",
    "1111101110100111",
    "1111101000011011",
    "1111100001110110",
    "1111011100000100",
    "1111011000000011",
    "1111010110010011",
    "1111010110111111",
    "1111011001110000",
    "1111011110000100",
    "1111100011001101",
    "1111101000011000",
    "1111101100101001",
    "1111101111000000",
    "1111101110101110",
    "1111101011011101",
    "1111100101100111",
    "1111011110010111",
    "1111010111010011",
    "1111010010001011",
    "1111010000001101",
    "1111010001111001",
    "1111010111000001",
    "1111011110110000",
    "1111101000001100",
    "1111110010011000",
    "1111111100011101",
    "1111111010011001",
    "1111110011001111",
    "1111101111000001",
    "1111101110101000",
    "1111110010100000",
    "1111111010001110",
    "1111111011011001",
    "1111110000011001",
    "1111100110111001",
    "1111100000111001",
    "1111011111111010",
    "1111100100101110",
    "1111101111011010",
    "1111111111001111",
    "1111101101011011",
    "1111011000111010",
    "1111000101101100",
    "1110110110000011",
    "1110101011100101",
    "1110100110111100",
    "1110100111111010",
    "1110101101101110",
    "1110110111011010",
    "1111000100000001",
    "1111010010101110",
    "1111100010011100",
    "1111110001101111",
    "1111111110111100",
    "1111110111101100",
    "1111110011100110",
    "1111110101010011",
    "1111111100001110",
    "1111111001010010",
    "1111101101110011",
    "1111100011111001",
    "1111011101111000",
    "1111011101001010",
    "1111100010000101",
    "1111101011111010",
    "1111111001000010",
    "1111111000101111",
    "1111101011110000",
    "1111100001111011",
    "1111011100101011",
    "1111011100101000",
    "1111100001100100",
    "1111101010011100",
    "1111110101100111",
    "1111111110111000",
    "1111110101000000",
    "1111101110010111",
    "1111101100000001",
    "1111101110011000",
    "1111110101010010",
    "1111111111111011",
    "1111110011001001",
    "1111100110000001",
    "1111011010111111",
    "1111010100001010",
    "1111010010111110",
    "1111010111110111",
    "1111100010000000",
    "1111101111101010",
    "1111111110100010",
    "1111110011011111",
    "1111101000001100",
    "1111100000100100",
    "1111011100111111",
    "1111011101010100",
    "1111100001000000",
    "1111100111011110",
    "1111101111111101",
    "1111111001101111",
    "1111111011111001",
    "1111110001110110",
    "1111101000111110",
    "1111100010000110",
    "1111011110001010",
    "1111011101111101",
    "1111100010000101",
    "1111101010101011",
    "1111110111001010",
    "1111111001111010",
    "1111101010101011",
    "1111011101010111",
    "1111010011111011",
    "1111001111011010",
    "1111010000000000",
    "1111010101000001",
    "1111011101010110",
    "1111100111110000",
    "1111110011000011",
    "1111111110000110",
    "1111111000001010",
    "1111110000110101",
    "1111101100110100",
    "1111101100101011",
    "1111110000011010",
    "1111110111001000",
    "1111111111010001",
    "1111111001001110",
    "1111110100011110",
    "1111110011111101",
    "1111111000011101",
    "1111111110001110",
    "1111110001010011",
    "1111100010011111",
    "1111010011111011",
    "1111000111100101",
    "1110111111000111",
    "1110111011101000",
    "1110111101101001",
    "1111000101000011",
    "1111010000111001",
    "1111011111100001",
    "1111101110100010",
    "1111111011010000",
    "1111111100101101",
    "1111111011000001",
    "1111111111111111",
    "1111110101100100",
    "1111101000001011",
    "1111011010111100",
    "1111010000110011",
    "1111001011110101",
    "1111001100111100",
    "1111010011101100",
    "1111011110110101",
    "1111101100010100",
    "1111111001111101",
    "1111111010010000",
    "1111110010000100",
    "1111101110100100",
    "1111110000011111",
    "1111111000001100",
    "1111111010100110",
    "1111101001000111",
    "1111010101011010",
    "1111000010001101",
    "1110110010010000",
    "1110100111101010",
    "1110100011011101",
    "1110100101010011",
    "1110101100000001",
    "1110110110000100",
    "1111000010100001",
    "1111010000111011",
    "1111100001001100",
    "1111110010110110",
    "1111111011010001",
    "1111101011001011",
    "1111011111000101",
    "1111011000111100",
    "1111011001110010",
    "1111100001010100",
    "1111101101111101",
    "1111111101001000",
    "1111110100000000",
    "1111101000000111",
    "1111100001000101",
    "1111011111111111",
    "1111100101000000",
    "1111101111100000",
    "1111111110001000",
    "1111110001000100",
    "1111100000010111",
    "1111010001111001",
    "1111000111011010",
    "1111000010000101",
    "1111000010100001",
    "1111001000110100",
    "1111010100011100",
    "1111100100010000",
    "1111110110011110",
    "1111110111001000",
    "1111100111001010",
    "1111011011101101",
    "1111010110001011",
    "1111010110110100",
    "1111011100101110",
    "1111100110000110",
    "1111110000101001",
    "1111111010001001",
    "1111111110111000",
    "1111111011000111",
    "1111111010010110",
    "1111111100000010",
    "1111111111101010",
    "1111111011001000",
    "1111110100110100",
    "1111101101111100",
    "1111100111010101",
    "1111100001111101",
    "1111011110101001",
    "1111011101111010",
    "1111011111101000",
    "1111100011010000",
    "1111101000000110",
    "1111101101100110",
    "1111110011101001",
    "1111111010100010",
    "1111111101010001",
    "1111110011101010",
    "1111101001000100",
    "1111011110110110",
    "1111010110111011",
    "1111010011010111",
    "1111010101100101",
    "1111011101101001",
    "1111101010010101",
    "1111111001001011",
    "1111111000100100",
    "1111101101011111",
    "1111100111010100",
    "1111100110101111",
    "1111101011100101",
    "1111110101001001",
    "1111111101011100",
    "1111101101010000",
    "1111011011010110",
    "1111001001001100",
    "1110111000100101",
    "1110101011011000",
    "1110100011010011",
    "1110100001011110",
    "1110100110000110",
    "1110110000101011",
    "1110111111111111",
    "1111010010001000",
    "1111100100110110",
    "1111110101101101",
    "1111111101011111",
    "1111110110010101",
    "1111110101011100",
    "1111111010011111",
    "1111111011101111",
    "1111101111000001",
    "1111100001001100",
    "1111010011111100",
    "1111001000101111",
    "1111000000110001",
    "1110111101000010",
    "1110111110010010",
    "1111000101001000",
    "1111010001100100",
    "1111100010110001",
    "1111110110111101",
    "1111110100010100",
    "1111100001101110",
    "1111010011010011",
    "1111001010001100",
    "1111000110100101",
    "1111001000000011",
    "1111001110001100",
    "1111011000110111",
    "1111101000000000",
    "1111111010111100",
    "1111101111110110",
    "1111011011000001",
    "1111001001100011",
    "1110111110011011",
    "1110111011110011",
    "1111000010101001",
    "1111010010010111",
    "1111101000111110",
    "1111111100101000",
    "1111100010000011",
    "1111001010100101",
    "1110111000101100",
    "1110101101101001",
    "1110101001100111",
    "1110101011110000",
    "1110110011000000",
    "1110111110101101",
    "1111001110100110",
    "1111100010100110",
    "1111111001110110",
    "1111101101011011",
    "1111010110010011",
    "1111000100001101",
    "1110111010001110",
    "1110111010000001",
    "1111000011001000",
    "1111010010110110",
    "1111100101001000",
    "1111110101100110",
    "1111111110111011",
    "1111111010001001",
    "1111111011110101",
    "1111111101011011",
    "1111110011101110",
    "1111101000101000",
    "1111011101001100",
    "1111010001110001",
    "1111000110100100",
    "1110111100000101",
    "1110110011101100",
    "1110101111010111",
    "1110110001011111",
    "1110111011111000",
    "1111001110110001",
    "1111101000001010",
    "1111111011100111",
    "1111100001001101",
    "1111001100101011",
    "1111000000101110",
    "1110111110011001",
    "1111000101001000",
    "1111010011001111",
    "1111100110010000",
    "1111111011011110",
    "1111101111110010",
    "1111011101111101",
    "1111010000111110",
    "1111001010000111",
    "1111001010001110",
    "1111010001111011",
    "1111100001011001",
    "1111110111111001",
    "1111101100101101",
    "1111010000000010",
    "1110110110010011",
    "1110100011100100",
    "1110011010101000",
    "1110011100100101",
    "1110101000101100",
    "1110111100101010",
    "1111010101010011",
    "1111101111001010",
    "1111111000110011",
    "1111100100111100",
    "1111010110101010",
    "1111001110101001",
    "1111001101010001",
    "1111010010110110",
    "1111011111011010",
    "1111110010000110",
    "1111110110111011",
    "1111011110110101",
    "1111001001001011",
    "1110111001010101",
    "1110110001110011",
    "1110110011110011",
    "1110111111000100",
    "1111010001111110",
    "1111101001110010",
    "1111111100110000",
    "1111100100101111",
    "1111010000011001",
    "1111000000110011",
    "1110110110001101",
    "1110110000001101",
    "1110101110010100",
    "1110110000010001",
    "1110110110001110",
    "1111000000100111",
    "1111001111110001",
    "1111100011010011",
    "1111111001101100",
    "1111101111110000",
    "1111011100100110",
    "1111010000000111",
    "1111001100011110",
    "1111010001111000",
    "1111011110011111",
    "1111101111001110",
    "1111111111010111",
    "1111110000000000",
    "1111100100010101",
    "1111011101000000",
    "1111011010001110",
    "1111011100000100",
    "1111100010111001",
    "1111101111001101",
    "1111111110111001",
    "1111101000011000",
    "1111001111010110",
    "1110110110110110",
    "1110100010001011",
    "1110010100000000",
    "1110001101110011",
    "1110001111101100",
    "1110011000101100",
    "1110100111001000",
    "1110111001010001",
    "1111001101101000",
    "1111100010111001",
    "1111111000000101",
    "1111110011111010",
    "1111100010011100",
    "1111010100110110",
    "1111001100011110",
    "1111001010001111",
    "1111001110011011",
    "1111011000011101",
    "1111100111000110",
    "1111111000101010",
    "1111110100100101",
    "1111100010010101",
    "1111010001111101",
    "1111000100101110",
    "1110111011100001",
    "1110110111000001",
    "1110110111010011",
    "1110111100000101",
    "1111000100101001",
    "1111001111111000",
    "1111011100100011",
    "1111101001011110",
    "1111110101101111",
    "1111111111001101",
    "1111110101111001",
    "1111101110101010",
    "1111101001111011",
    "1111100111111100",
    "1111101000101111",
    "1111101011111111",
    "1111110000111011",
    "1111110110100101",
    "1111111011111011",
    "1111111111110000",
    "1111111101000010",
    "1111111100000010",
    "1111111100101100",
    "1111111110110100",
    "1111111101110010",
    "1111111001011110",
    "1111110100011110",
    "1111101111001010",
    "1111101001111111",
    "1111100101101001",
    "1111100010101111",
    "1111100010000010",
    "1111100100000101",
    "1111101001010011",
    "1111110001110000",
    "1111111101000001",
    "1111110101110110",
    "1111101000011011",
    "1111011100100001",
    "1111010011111000",
    "1111001111110001",
    "1111010000110000",
    "1111010110100000",
    "1111100000000010",
    "1111101011110010",
    "1111111000000110",
    "1111111100101100",
    "1111110100000011",
    "1111101110110001",
    "1111101101000101",
    "1111101110101000",
    "1111110010101011",
    "1111111000010100",
    "1111111110101100",
    "1111111011000001",
    "1111110101101000",
    "1111110001110010",
    "1111110000000110",
    "1111110000111111",
    "1111110100101110",
    "1111111011010011",
    "1111111011110001",
    "1111110001011111",
    "1111100111001010",
    "1111011110001101",
    "1111010111111110",
    "1111010101001101",
    "1111010110000011",
    "1111011001111100",
    "1111011111110000",
    "1111100110011010",
    "1111101100111100",
    "1111110010110111",
    "1111111000000111",
    "1111111100111110",
    "1111111110001101",
    "1111111001011011",
    "1111110100110110",
    "1111110001000111",
    "1111101111000010",
    "1111101111010110",
    "1111110010100011",
    "1111111000100110",
    "1111111111000100",
    "1111110101100010",
    "1111101100000110",
    "1111100100000101",
    "1111011110011011",
    "1111011011101011",
    "1111011011110010",
    "1111011110001111",
    "1111100010001010",
    "1111100110101000",
    "1111101010111010",
    "1111101110101000",
    "1111110001101010",
    "1111110100010000",
    "1111110110101000",
    "1111111000111011",
    "1111111011000100",
    "1111111100110101",
    "1111111101111010",
    "1111111110001101",
    "1111111101111000",
    "1111111101011011",
    "1111111101100000",
    "1111111110101100",
    "1111111110101010",
    "1111111010110110",
    "1111110110011100",
    "1111110010011011",
    "1111101111101111",
    "1111101110111110",
    "1111110000001000",
    "1111110010100110",
    "1111110101011110",
    "1111110111110110",
    "1111111001001011",
    "1111111001011001",
    "1111111001000100",
    "1111111001000010",
    "1111111010010010",
    "1111111101100011",
    "1111111100110100",
    "1111110101000100",
    "1111101011111001",
    "1111100010011010",
    "1111011001111100",
    "1111010011101100",
    "1111010000100111",
    "1111010001001010",
    "1111010101011011",
    "1111011101001100",
    "1111100111111110",
    "1111110101001011",
    "1111111100000110",
    "1111101101001101",
    "1111011111101000",
    "1111010100110001",
    "1111001101110010",
    "1111001011000110",
    "1111001100011011",
    "1111010000111000",
    "1111010111011101",
    "1111011111011001",
    "1111101000010101",
    "1111110010011011",
    "1111111101110010",
    "1111110101110101",
    "1111101001011101",
    "1111011110100011",
    "1111010110101111",
    "1111010011001010",
    "1111010100000001",
    "1111011000100111",
    "1111011111011010",
    "1111100110110001",
    "1111101101010001",
    "1111110010001101",
    "1111110101010101",
    "1111110110110010",
    "1111110110110001",
    "1111110101011001",
    "1111110010101111",
    "1111101111000011",
    "1111101010101110",
    "1111100110011110",
    "1111100011000101",
    "1111100001010000",
    "1111100001011001",
    "1111100011011010",
    "1111100111000101",
    "1111101011111100",
    "1111110001011001",
    "1111110110110001",
    "1111111011010100",
    "1111111110010010",
    "1111111111010000",
    "1111111110001110",
    "1111111011110011",
    "1111111001000101",
    "1111110111011000",
    "1111110111101111",
    "1111111010110011",
    "1111111111100101",
    "1111111000010010",
    "1111110000100111",
    "1111101010001010",
    "1111100110001110",
    "1111100101101110",
    "1111101000110000",
    "1111101110111101",
    "1111110111010101",
    "1111111111011010",
    "1111110110110110",
    "1111110000011010",
    "1111101101001111",
    "1111101101111001",
    "1111110010001111",
    "1111111001011110",
    "1111111101101110",
    "1111110100110011",
    "1111101101000000",
    "1111100111001001",
    "1111100011100100",
    "1111100010001111",
    "1111100010110011",
    "1111100100111011",
    "1111101000010000",
    "1111101100101010",
    "1111110010000110",
    "1111111000011111",
    "1111111111100100",
    "1111111001001101",
    "1111110010100111",
    "1111101101010011",
    "1111101001101101",
    "1111101000000000",
    "1111101000000100",
    "1111101001100011",
    "1111101100000000",
    "1111101110111000",
    "1111110001100110",
    "1111110011101001",
    "1111110100101011",
    "1111110100100000",
    "1111110011001001",
    "1111110000101111",
    "1111101101100000",
    "1111101001100111",
    "1111100101001110",
    "1111100000101001",
    "1111011100001111",
    "1111011000101100",
    "1111010110110111",
    "1111010111110100",
    "1111011100100110",
    "1111100110000011",
    "1111110100010111",
    "1111111000111100",
    "1111100011011111",
    "1111001101010100",
    "1110111000101100",
    "1110100111100000",
    "1110011011000111",
    "1110010011111001",
    "1110010001011110",
    "1110010010110011",
    "1110010110100010",
    "1110011011011001",
    "1110100000010100",
    "1110100100100100",
    "1110100111101111",
    "1110101001111010",
    "1110101011010110",
    "1110101100010100",
    "1110101101001001",
    "1110101101111011",
    "1110101110101110",
    "1110101111011110",
    "1110110000000000",
    "1110110000011100",
    "1110110001101100",
    "1110110110000000",
    "1110111111101001",
    "1111001111011111",
    "1111100100001011",
    "1111111010100000",
    "1111110001001100",
    "1111100001110001",
    "1111011000001001",
    "1111010010110011",
    "1111001110101001",
    "1111001000101010",
    "1110111111010110",
    "1110110011001011",
    "1110100110010000",
    "1110011011001010",
    "1110010100001011",
    "1110010010010010",
    "1110010100111100",
    "1110011010100011",
    "1110100001000010",
    "1110100110101100",
    "1110101010100010",
    "1110101100101011",
    "1110101110000101",
    "1110110000001100",
    "1110110100010010",
    "1110111011000110",
    "1111000100011101",
    "1111001111000000",
    "1111011000011010",
    "1111011110010100",
    "1111011111001101",
    "1111011011000110",
    "1111010011011000",
    "1111001010100010",
    "1111000010111101",
    "1110111110011001",
    "1110111101100110",
    "1111000000001010",
    "1111000101000001",
    "1111001010111000",
    "1111010000110001",
    "1111010110000011",
    "1111011010100011",
    "1111011110010001",
    "1111100001001111",
    "1111100011010011",
    "1111100100011101",
    "1111100100110100",
    "1111100100110111",
    "1111100101011010",
    "1111100111000011",
    "1111101010000110",
    "1111101110010011",
    "1111110010111100",
    "1111110111001100",
    "1111111010010110",
    "1111111011111010",
    "1111111011110000",
    "1111111001111101",
    "1111110110110011",
    "1111110010100110",
    "1111101101100101",
    "1111101000000100",
    "1111100010011101",
    "1111011101011001",
    "1111011001100000",
    "1111010111010101",
    "1111010111000110",
    "1111011000110010",
    "1111011011111101",
    "1111100000000011",
    "1111100100010011",
    "1111101000000101",
    "1111101010110111",
    "1111101100010111",
    "1111101100100001",
    "1111101011100101",
    "1111101001111010",
    "1111101000000010",
    "1111100110011110",
    "1111100101101001",
    "1111100101110110",
    "1111100111010111",
    "1111101010001100",
    "1111101110010011",
    "1111110011100010",
    "1111111001101101",
    "1111111111011000",
    "1111111000000100",
    "1111110000101011",
    "1111101001100101",
    "1111100011010000",
    "1111011110000010",
    "1111011010001011",
    "1111010111100111",
    "1111010110001001",
    "1111010101011011",
    "1111010101001001",
    "1111010101000110",
    "1111010101001011",
    "1111010101011111",
    "1111010110000011",
    "1111010110110001",
    "1111010111010001",
    "1111010111000011",
    "1111010101011011",
    "1111010010000010",
    "1111001100101101",
    "1111000101101111",
    "1110111101110010",
    "1110110101101110",
    "1110101110011111",
    "1110101000111100",
    "1110100101100111",
    "1110100100101010",
    "1110100101111100",
    "1110101001000010",
    "1110101101011110",
    "1110110010110001",
    "1110111000100111",
    "1110111110101110",
    "1111000100110001",
    "1111001010011000",
    "1111001111001010",
    "1111010010110110",
    "1111010101010111",
    "1111010110110100",
    "1111010111101000",
    "1111011000001110",
    "1111011000111111",
    "1111011010001001",
    "1111011011100011",
    "1111011100110010",
    "1111011101010100",
    "1111011100100001",
    "1111011001111001",
    "1111010101001000",
    "1111001110001100",
    "1111000101100100",
    "1110111100001100",
    "1110110011100100",
    "1110101101001111",
    "1110101010100010",
    "1110101100000101",
    "1110110001110001",
    "1110111010101011",
    "1111000101100111",
    "1111010001010101",
    "1111011100111101",
    "1111100111110001",
    "1111110001001001",
    "1111111000011011",
    "1111111101000000",
    "1111111110100010",
    "1111111100111100",
    "1111111000101110",
    "1111110010101100",
    "1111101011110100",
    "1111100100110110",
    "1111011110000101",
    "1111010111101000",
    "1111010001011001",
    "1111001011011011",
    "1111000110001000",
    "1111000010001101",
    "1111000000001111",
    "1111000000100001",
    "1111000010110011",
    "1111000110010011",
    "1111001010000110",
    "1111001101010100",
    "1111001111100110",
    "1111010001000010",
    "1111010001111110",
    "1111010010110100",
    "1111010011110100",
    "1111010100111100",
    "1111010110000011",
    "1111010111000011",
    "1111011000001000",
    "1111011001101011",
    "1111011100001111",
    "1111011111111111",
    "1111100100101111",
    "1111101001111010",
    "1111101110100101",
    "1111110001111110",
    "1111110011100110",
    "1111110011011011",
    "1111110001111000",
    "1111101111101011",
    "1111101101101001",
    "1111101100100100",
    "1111101101000100",
    "1111101111100010",
    "1111110100000010",
    "1111111010010001",
    "1111111110100001",
    "1111110111100010",
    "1111110001111111",
    "1111101110111101",
    "1111101111000010",
    "1111110010001111",
    "1111111000000000",
    "1111111111010110",
    "1111111000111010",
    "1111110010000011",
    "1111101101000000",
    "1111101010100010",
    "1111101010111110",
    "1111101110010011",
    "1111110100001011",
    "1111111011111110",
    "1111111010111001",
    "1111110001000111",
    "1111100111001010",
    "1111011101100110",
    "1111010101000001",
    "1111001110000010",
    "1111001000111110",
    "1111000110000000",
    "1111000101000011",
    "1111000101111100",
    "1111001000011010",
    "1111001100010011",
    "1111010001010010",
    "1111010110111110",
    "1111011100110000",
    "1111100001110100",
    "1111100101100111",
    "1111100111110011",
    "1111101000011111",
    "1111101000001100",
    "1111100111100101",
    "1111100111001110",
    "1111100111100010",
    "1111101000101011",
    "1111101010100101",
    "1111101101001010",
    "1111110000010010",
    "1111110011111101",
    "1111111000010001",
    "1111111101010001",
    "1111111101000111",
    "1111110111011101",
    "1111110010100100",
    "1111101111011111",
    "1111101111001000",
    "1111110001111010",
    "1111110111010111",
    "1111111110010101",
    "1111111010101001",
    "1111110100111001",
    "1111110001000010",
    "1111101110111011",
    "1111101101110000",
    "1111101100100000",
    "1111101010010110",
    "1111100110110111",
    "1111100010000010",
    "1111011100000001",
    "1111010101001011",
    "1111001101111000",
    "1111000110100000",
    "1110111111011110",
    "1110111001010011",
    "1110110101000011",
    "1110110100001010",
    "1110111000000001",
    "1111000001011100",
    "1111001111111101",
    "1111100001101011",
    "1111110011100101",
    "1111111101011011",
    "1111110011110110",
    "1111110000100010",
    "1111110010110000",
    "1111111000111010",
    "1111111110011000",
    "1111110011001101",
    "1111100011111001",
    "1111001110100100",
    "1110110011000110",
    "1110010011111110",
    "1101110101111110",
    "1101011110100100",
    "1101010001110110",
    "1101010001000000",
    "1101011001100111",
    "1101100110110100",
    "1101110011011111",
    "1101111100000111",
    "1101111111101100",
    "1101111111010010",
    "1101111100111111",
    "1101111010101010",
    "1101111001011011",
    "1101111001010000",
    "1101111001011001",
    "1101111001001001",
    "1101111000000110",
    "1101110110100000",
    "1101110100111011",
    "1101110011111110",
    "1101110011111100",
    "1101110101000101",
    "1101110111101111",
    "1101111101011001",
    "1110001000101101",
    "1110011100010110",
    "1110111001101010",
    "1111011111010111",
    "1111110110110101",
    "1111001111000010",
    "1110101111001000",
    "1110011011001110",
    "1110010011110011",
    "1110010110001101",
    "1110011110000100",
    "1110100110111111",
    "1110101110001100",
    "1110110010110110",
    "1110110101011101",
    "1110110111001101",
    "1110111000110111",
    "1110111010100101",
    "1110111100000010",
    "1110111100111100",
    "1110111101000111",
    "1110111100101110",
    "1110111100000001",
    "1110111011000001",
    "1110111001100010",
    "1110110111001001",
    "1110110011111000",
    "1110110000000101",
    "1110101100100110",
    "1110101010011000",
    "1110101010000100",
    "1110101100000101",
    "1110110001001111",
    "1110111011101010",
    "1111001110000000",
    "1111101001101100",
    "1111110010011110",
    "1111001011000010",
    "1110100110011000",
    "1110001010111100",
    "1101111101001100",
    "1101111101111111",
    "1110001010010110",
    "1110011101001001",
    "1110110001001010",
    "1111000011001011",
    "1111010010100111",
    "1111100000100110",
    "1111101110110001",
    "1111111101111101",
    "1111110010100110",
    "1111100100111110",
    "1111011011011001",
    "1111010111010101",
    "1111011000011101",
    "1111011101000010",
    "1111100010101001",
    "1111100111100010",
    "1111101011000000",
    "1111101101010110",
    "1111101111001110",
    "1111110001001000",
    "1111110010111010",
    "1111110011110010",
    "1111110010100000",
    "1111101101111111",
    "1111100101110100",
    "1111011010011101",
    "1111001101001111",
    "1111000000000010",
    "1110110100101010",
    "1110101100100101",
    "1110101000101101",
    "1110101001010011",
    "1110101101111111",
    "1110110101110100",
    "1110111111100011",
    "1111001001101111",
    "1111010011001010",
    "1111011011000010",
    "1111100001001010",
    "1111100101111001",
    "1111101001110010",
    "1111101101011100",
    "1111110001011010",
    "1111110110001100",
    "1111111100010111",
    "1111111011100111",
    "1111110001111001",
    "1111100111000101",
    "1111011100100000",
    "1111010011101111",
    "1111001110010110",
    "1111001101010100",
    "1111010000111000",
    "1111011000010000",
    "1111100010000010",
    "1111101100011110",
    "1111110110000011",
    "1111111101101101",
    "1111111101000110",
    "1111111010100000",
    "1111111010001100",
    "1111111011110011",
    "1111111111000001",
    "1111111100010000",
    "1111110110001001",
    "1111101110100011",
    "1111100101101111",
    "1111011100010001",
    "1111010011000001",
    "1111001011000100",
    "1111000101010011",
    "1111000010010010",
    "1111000001111110",
    "1111000011111110",
    "1111000111101100",
    "1111001100101000",
    "1111010010100111",
    "1111011001101101",
    "1111100001111000",
    "1111101010101011",
    "1111110011000111",
    "1111111001110011",
    "1111111101011111",
    "1111111101100111",
    "1111111010100000",
    "1111110101011101",
    "1111110000010110",
    "1111101100111101",
    "1111101100011100",
    "1111101111000111",
    "1111110100011100",
    "1111111011011001",
    "1111111101000011",
    "1111110101110101",
    "1111101111011010",
    "1111101010000000",
    "1111100101101100",
    "1111100010011010",
    "1111100000001000",
    "1111011110110110",
    "1111011110011110",
    "1111011110110101",
    "1111011111101001",
    "1111100000110000",
    "1111100010001000",
    "1111100011111110",
    "1111100110100001",
    "1111101010000010",
    "1111101110100101",
    "1111110011111101",
    "1111111001110110",
    "1111111111111001",
    "1111111010001001",
    "1111110100100000",
    "1111101111010111",
    "1111101010111100",
    "1111100111100101",
    "1111100101101010",
    "1111100101011000",
    "1111100110110001",
    "1111101001011111",
    "1111101101000010",
    "1111110000101101",
    "1111110011110000",
    "1111110101011111",
    "1111110101011101",
    "1111110011011111",
    "1111101111111001",
    "1111101011010110",
    "1111100110101101",
    "1111100010110110",
    "1111100000010111",
    "1111011111100100",
    "1111100000011001",
    "1111100010100111",
    "1111100101110010",
    "1111101001100110",
    "1111101101101010",
    "1111110001101111",
    "1111110101101001",
    "1111111001001010",
    "1111111100001011",
    "1111111110101001",
    "1111111111011001",
    "1111111110000100",
    "1111111101011000",
    "1111111101010110",
    "1111111101110111",
    "1111111110110010",
    "1111111111111001",
    "1111111111000111",
    "1111111110101111",
    "1111111111011111",
    "1111111110001000",
    "1111111001110000",
    "1111110011001111",
    "1111101010110100",
    "1111100001000011",
    "1111010110110111",
    "1111001101001010",
    "1111000100100111",
    "1110111101101110",
    "1110111000101101",
    "1110110101101010",
    "1110110100101100",
    "1110110101101111",
    "1110111000101000",
    "1110111100111101",
    "1111000010000011",
    "1111000111001001",
    "1111001011010110",
    "1111001110000101",
    "1111001111001010",
    "1111001111000100",
    "1111001110110000",
    "1111001111010010",
    "1111010001011010",
    "1111010101010101",
    "1111011010100101",
    "1111100000010100",
    "1111100101101001",
    "1111101001110011",
    "1111101100011001",
    "1111101101001111",
    "1111101100010010",
    "1111101001101000",
    "1111100101011010",
    "1111011111111010",
    "1111011001010110",
    "1111010001111000",
    "1111001001101011",
    "1111000001010111",
    "1110111010000001",
    "1110110101001000",
    "1110110100001000",
    "1110110111110111",
    "1111000000000111",
    "1111001011100110",
    "1111011000011010",
    "1111100100101110",
    "1111101111011100",
    "1111111000011010",
    "1111111111111110",
    "1111111001010110",
    "1111110011100110",
    "1111101111001110",
    "1111101100111100",
    "1111101101010111",
    "1111110000100011",
    "1111110101110100",
    "1111111011111010",
    "1111111110011111",
    "1111111010011111",
    "1111111000011100",
    "1111111000001011",
    "1111111001000010",
    "1111111010010000",
    "1111111011001101",
    "1111111011011111",
    "1111111011000011",
    "1111111010000001",
    "1111111000100101",
    "1111110110110101",
    "1111110100101011",
    "1111110001111011",
    "1111101110011010",
    "1111101010010101",
    "1111100110001011",
    "1111100010101011",
    "1111100000011001",
    "1111011111100100",
    "1111011111110001",
    "1111100000000000",
    "1111011110111111",
    "1111011011101000",
    "1111010101100010",
    "1111001101001010",
    "1111000100000110",
    "1110111100011100",
    "1110111000011110",
    "1110111001110010",
    "1111000001000010",
    "1111001101100110",
    "1111011101110101",
    "1111101111011011",
    "1111111111111100",
    "1111110010010010",
    "1111101000101111",
    "1111100011110100",
    "1111100011101010",
    "1111101000011100",
    "1111110010100000",
    "1111111110001010",
    "1111101010011110",
    "1111010100100010",
    "1110111111011001",
    "1110101110011011",
    "1110100100010010",
    "1110100010011010",
    "1110101000101010",
    "1110110101110001",
    "1111001000000100",
    "1111011110000101",
    "1111110110010111",
    "1111110000101101",
    "1111011001010001",
    "1111000101011010",
    "1110110111000001",
    "1110101111000111",
    "1110101101100110",
    "1110110001001000",
    "1110110111100011",
    "1110111110100011",
    "1111000100011010",
    "1111001000010101",
    "1111001010001111",
    "1111001010101000",
    "1111001001111010",
    "1111001000010000",
    "1111000101101001",
    "1111000001111110",
    "1110111101001111",
    "1110110111101101",
    "1110110001110011",
    "1110101100000101",
    "1110100111000100",
    "1110100011001101",
    "1110100000111001",
    "1110100000011111",
    "1110100010010100",
    "1110100110011011",
    "1110101100101110",
    "1110110100111001",
    "1110111110011110",
    "1111001010010100",
    "1111011011001001",
    "1111110011100001",
    "1111101011111110",
    "1111000110001001",
    "1110100000100100",
    "1110000001101100",
    "1101101110110110",
    "1101101010010001",
    "1101110001110001",
    "1101111111111011",
    "1110001110100110",
    "1110011001001001",
    "1110011101110111",
    "1110011101100110",
    "1110011010100011",
    "1110010111000110",
    "1110010100110110",
    "1110010011111011",
    "1110010011100110",
    "1110010010111110",
    "1110010001100111",
    "1110001111110011",
    "1110001110011011",
    "1110001110001100",
    "1110001111010100",
    "1110010001100001",
    "1110010100101010",
    "1110011000111010",
    "1110011110011110",
    "1110100101100000",
    "1110101110000100",
    "1110111000100010",
    "1111000110101010",
    "1111011010110111",
    "1111110110010111",
    "1111100111111001",
    "1111000011110100",
    "1110100011000001",
    "1110001011000001",
    "1101111111100001",
    "1110000000110000",
    "1110001011001110",
    "1110011001101111",
    "1110100111001101",
    "1110110000100100",
    "1110110101100101",
    "1110110111111100",
    "1110111010011101",
    "1110111111100001",
    "1111000111111010",
    "1111010010110001",
    "1111011110010001",
    "1111101000100101",
    "1111110000100111",
    "1111110110010111",
    "1111111010001110",
    "1111111100100001",
    "1111111101011011",
    "1111111100111111",
    "1111111011011101",
    "1111111001001001",
    "1111110110101110",
    "1111110101000110",
    "1111110101001101",
    "1111110111100111",
    "1111111100011000",
    "1111111100111101",
    "1111110101011110",
    "1111101110010101",
    "1111101000110011",
    "1111100101111110",
    "1111100110011101",
    "1111101010011000",
    "1111110001010001",
    "1111111010001000",
    "1111111100010100",
    "1111110011101011",
    "1111101101001001",
    "1111101001001111",
    "1111100111101111",
    "1111100111110100",
    "1111101000100011",
    "1111101001001101",
    "1111101001010010",
    "1111101000010100",
    "1111100101111100",
    "1111100001110100",
    "1111011011111101",
    "1111010100110001",
    "1111001101001010",
    "1111000110010000",
    "1111000001001111",
    "1110111110111000",
    "1110111111011100",
    "1111000010010000",
    "1111000110010000",
    "1111001010000111",
    "1111001100101110",
    "1111001101011110",
    "1111001100001010",
    "1111001001001100",
    "1111000101010101",
    "1111000001010101",
    "1110111101110011",
    "1110111010111101",
    "1110111000110010",
    "1110110111000110",
    "1110110101101010",
    "1110110100011010",
    "1110110011010000",
    "1110110010010100",
    "1110110001101100",
    "1110110001100111",
    "1110110010010010",
    "1110110011110011",
    "1110110110001000",
    "1110111000111111",
    "1110111011111101",
    "1110111110100001",
    "1111000000010001",
    "1111000001000101",
    "1111000001000111",
    "1111000000101100",
    "1111000000011001",
    "1111000000110101",
    "1111000010100100",
    "1111000101111001",
    "1111001010110101",
    "1111010001001100",
    "1111011000101010",
    "1111100001000000",
    "1111101001111101",
    "1111110011001100",
    "1111111100010101",
    "1111111011000100",
    "1111110011011111",
    "1111101101001000",
    "1111101000001000",
    "1111100100100010",
    "1111100010011100",
    "1111100010000110",
    "1111100011101010",
    "1111100110111011",
    "1111101011010100",
    "1111101111111110",
    "1111110100001100",
    "1111110111101101",
    "1111111010111000",
    "1111111110011001",
    "1111111101000010",
    "1111110111010001",
    "1111110000101001",
    "1111101001111111",
    "1111100100010000",
    "1111100000000011",
    "1111011101101101",
    "1111011101000101",
    "1111011101111111",
    "1111100000010001",
    "1111100011110011",
    "1111101000100100",
    "1111101110011000",
    "1111110100111011",
    "1111111011100111",
    "1111111110010010",
    "1111111001101111",
    "1111110111011110",
    "1111111000000011",
    "1111111011100100",
    "1111111110011000",
    "1111110110110110",
    "1111101111000001",
    "1111100111111100",
    "1111100010001000",
    "1111011101100000",
    "1111011001100101",
    "1111010101110111",
    "1111010010001000",
    "1111001110101011",
    "1111001100010100",
    "1111001100000010",
    "1111001110100011",
    "1111010011111001",
    "1111011011010100",
    "1111100011100111",
    "1111101011011011",
    "1111110001100110",
    "1111110101011110",
    "1111110111000001",
    "1111110110110001",
    "1111110101100111",
    "1111110100100101",
    "1111110100011111",
    "1111110101110010",
    "1111111000011110",
    "1111111100001001",
    "1111111111110010",
    "1111111011111010",
    "1111111000011000",
    "1111110101000111",
    "1111110001111011",
    "1111101110110100",
    "1111101100000110",
    "1111101010001111",
    "1111101001101100",
    "1111101010101010",
    "1111101100110101",
    "1111101111100000",
    "1111110001101000",
    "1111110010010010",
    "1111110001000100",
    "1111101110010010",
    "1111101010111001",
    "1111101000000101",
    "1111100110101110",
    "1111100111000000",
    "1111101000011110",
    "1111101010011001",
    "1111101100001100",
    "1111101101101110",
    "1111101111010001",
    "1111110001000111",
    "1111110011001111",
    "1111110101001001",
    "1111110110001001",
    "1111110101100010",
    "1111110011000101",
    "1111101111000111",
    "1111101010011011",
    "1111100110001000",
    "1111100011011010",
    "1111100011000110",
    "1111100101011000",
    "1111101001101100",
    "1111101110111101",
    "1111110011111011",
    "1111110111100000",
    "1111111001001000",
    "1111111000111110",
    "1111110111111111",
    "1111110111100001",
    "1111111000110010",
    "1111111100011100",
    "1111111101101100",
    "1111110110100111",
    "1111101111101011",
    "1111101010010001",
    "1111100111001010",
    "1111100110011010",
    "1111100111100100",
    "1111101010001000",
    "1111101101111000",
    "1111110010111000",
    "1111111001000110",
    "1111111111110110",
    "1111111001000001",
    "1111110011101110",
    "1111110001010011",
    "1111110010101100",
    "1111110111111111",
    "1111111111110000",
    "1111110110100101",
    "1111101110111001",
    "1111101011000011",
    "1111101100110010",
    "1111110100101100",
    "1111111101101100",
    "1111101011111011",
    "1111010111111100",
    "1111000011100010",
    "1110110000010100",
    "1110011111011111",
    "1110010010010000",
    "1110001001110000",
    "1110000111001000",
    "1110001011010001",
    "1110010110010110",
    "1110100111100011",
    "1110111100110000",
    "1111010010111011",
    "1111100110111001",
    "1111110110001011",
    "1111111111100111",
    "1111111100011011",
    "1111111100100100",
    "1111111110111111",
    "1111111101101110",
    "1111111010001001",
    "1111110101111011",
    "1111110000000000",
    "1111100111010001",
    "1111011011000100",
    "1111001011110010",
    "1110111010111101",
    "1110101011000010",
    "1110011110101000",
    "1110010111101100",
    "1110010111000011",
    "1110011100001010",
    "1110100101100010",
    "1110110001101011",
    "1110111111110000",
    "1111010000000111",
    "1111100011100100",
    "1111111010011000",
    "1111101100110101",
    "1111010101001000",
    "1111000010010010",
    "1110110111100000",
    "1110110110001001",
    "1110111101000000",
    "1111001000101111",
    "1111010101000101",
    "1111011110011011",
    "1111100010111011",
    "1111100010101110",
    "1111011111001111",
    "1111011010010110",
    "1111010101100000",
    "1111010001011001",
    "1111001101110111",
    "1111001010011000",
    "1111000110011111",
    "1111000010001000",
    "1110111101101001",
    "1110111001101000",
    "1110110110100000",
    "1110110100101100",
    "1110110100010111",
    "1110110101101100",
    "1110111000110010",
    "1110111101101001",
    "1111000100001011",
    "1111001100001100",
    "1111010110011010",
    "1111100100111110",
    "1111111010000100",
    "1111101001011110",
    "1111000111100000",
    "1110100100100000",
    "1110000110000110",
    "1101110001010010",
    "1101101000110010",
    "1101101011100011",
    "1101110101011010",
    "1110000000111110",
    "1110001001101010",
    "1110001101001110",
    "1110001011111100",
    "1110000111110001",
    "1110000011010101",
    "1110000000101001",
    "1110000000010100",
    "1110000001111011",
    "1110000100011101",
    "1110000111000011",
    "1110001001011001",
    "1110001011101101",
    "1110001110000101",
    "1110010000011010",
    "1110010010001010",
    "1110010010111001",
    "1110010010101001",
    "1110010001111000",
    "1110010001011010",
    "1110010011001111",
    "1110011010110101",
    "1110101011110111",
    "1111000111111110",
    "1111101101011000",
    "1111101001000101",
    "1111000010101001",
    "1110100110000000",
    "1110010111100000",
    "1110010111010000",
    "1110100001010000",
    "1110101111111010",
    "1110111101110111",
    "1111000111111110",
    "1111001101110000",
    "1111010000011100",
    "1111010010000101",
    "1111010100011111",
    "1111011000010011",
    "1111011101000101",
    "1111100001111101",
    "1111100101111100",
    "1111101000101111",
    "1111101010100101",
    "1111101011111111",
    "1111101101001111",
    "1111101110010110",
    "1111101111011001",
    "1111110000100100",
    "1111110001111111",
    "1111110011101000",
    "1111110101100100",
    "1111111000001000",
    "1111111100000010",
    "1111111101111010",
    "1111110101011010",
    "1111101010110011",
    "1111011111001010",
    "1111010100010011",
    "1111001100000100",
    "1111000111111010",
    "1111001000011011",
    "1111001101010010",
    "1111010101100010",
    "1111011111101011",
    "1111101010000010",
    "1111110011001011",
    "1111111010001110",
    "1111111111000100",
    "1111111101101110",
    "1111111011001111",
    "1111111000011100",
    "1111110100100110",
    "1111101111010000",
    "1111101000011111",
    "1111100000110001",
    "1111011000110111",
    "1111010001101100",
    "1111001100000101",
    "1111001000100111",
    "1111000111101010",
    "1111001001011011",
    "1111001101110011",
    "1111010100001011",
    "1111011011100110",
    "1111100010110110",
    "1111101000110000",
    "1111101100011111",
    "1111101101101110",
    "1111101100101011",
    "1111101001111111",
    "1111100110010010",
    "1111100001111001",
    "1111011101000101",
    "1111010111110001",
    "1111010001111000",
    "1111001011011001",
    "1111000100100100",
    "1110111101111011",
    "1110111000010000",
    "1110110100010111",
    "1110110010101111",
    "1110110011101110",
    "1110110111001011",
    "1110111100101110",
    "1111000011101010",
    "1111001011000010",
    "1111010001110001",
    "1111010110101100",
    "1111011000111100",
    "1111011000000100",
    "1111010100011100",
    "1111001111000010",
    "1111001001011101",
    "1111000101010101",
    "1111000100000011",
    "1111000110010011",
    "1111001100000100",
    "1111010100101110",
    "1111011111001101",
    "1111101010010110",
    "1111110100111100",
    "1111111110001001",
    "1111111010011101",
    "1111110101000101",
    "1111110001100110",
    "1111101111110101",
    "1111101111110000",
    "1111110001011011",
    "1111110100110011",
    "1111111001011110",
    "1111111110011001",
    "1111111101101100",
    "1111111100000101",
    "1111111101010001",
    "1111111111001100",
    "1111111010101001",
    "1111110110110001",
    "1111110101000000",
    "1111110110000001",
    "1111111001011000",
    "1111111101111110",
    "1111111101010111",
    "1111111001011011",
    "1111110110001011",
    "1111110011001000",
    "1111101111101100",
    "1111101011101010",
    "1111100111011010",
    "1111100011101010",
    "1111100001001010",
    "1111100000001101",
    "1111100000100111",
    "1111100001101110",
    "1111100010110001",
    "1111100011000110",
    "1111100010011100",
    "1111100000110110",
    "1111011110110101",
    "1111011101001001",
    "1111011100011110",
    "1111011101001111",
    "1111011111000111",
    "1111100001001111",
    "1111100010011100",
    "1111100001111011",
    "1111011111101011",
    "1111011100100011",
    "1111011001110111",
    "1111011000111010",
    "1111011010010011",
    "1111011101101101",
    "1111100010001011",
    "1111100110100001",
    "1111101001101101",
    "1111101011010111",
    "1111101011101110",
    "1111101011011101",
    "1111101011011011",
    "1111101100001110",
    "1111101110001000",
    "1111110000111111",
    "1111110100011100",
    "1111111000000011",
    "1111111011100011",
    "1111111110111011",
    "1111111101011100",
    "1111111001000101",
    "1111110011100001",
    "1111101100101110",
    "1111100101001101",
    "1111011101111111",
    "1111011000001001",
    "1111010100100010",
    "1111010011010010",
    "1111010011111001",
    "1111010101100000",
    "1111010111100000",
    "1111011001101011",
    "1111011100010100",
    "1111011111110101",
    "1111100100001011",
    "1111101000111100",
    "1111101101010001",
    "1111110000010001",
    "1111110001100011",
    "1111110001010110",
    "1111110000011110",
    "1111101111111110",
    "1111110000110001",
    "1111110011010011",
    "1111110111001111",
    "1111111011101010",
    "1111111111001111",
    "1111111111010011",
    "1111111110111001",
    "1111111001011100",
    "1111110000100001",
    "1111100101001011",
    "1111011001000001",
    "1111001101111111",
    "1111000101101001",
    "1111000001000111",
    "1111000000110101",
    "1111000100100100",
    "1111001011110010",
    "1111010101111110",
    "1111100010111110",
    "1111110010101101",
    "1111111011010110",
    "1111101000101011",
    "1111010111011010",
    "1111001010000110",
    "1111000010111110",
    "1111000011001000",
    "1111001010001001",
    "1111010110000001",
    "1111100011111001",
    "1111110001000101",
    "1111111011111000",
    "1111111100010000",
    "1111110111011001",
    "1111110101100110",
    "1111110111011000",
    "1111111101001111",
    "1111111001000011",
    "1111101100111001",
    "1111100000101011",
    "1111010111001000",
    "1111010010011100",
    "1111010011101010",
    "1111011010101011",
    "1111100110100111",
    "1111110110000000",
    "1111111000101111",
    "1111100111100101",
    "1111011000100000",
    "1111001101001111",
    "1111000110110100",
    "1111000101010000",
    "1111000111100111",
    "1111001100101010",
    "1111010011010000",
    "1111011010100110",
    "1111100010001000",
    "1111101001011011",
    "1111110000000001",
    "1111110101011101",
    "1111111001010000",
    "1111111011001010",
    "1111111011010100",
    "1111111010010101",
    "1111111001000001",
    "1111111000001001",
    "1111111000000110",
    "1111111000100110",
    "1111111000111000",
    "1111110111110111",
    "1111110100100100",
    "1111101110011001",
    "1111100101011000",
    "1111011010010011",
    "1111001110100011",
    "1111000011111100",
    "1110111100010100",
    "1110111001000110",
    "1110111011000111",
    "1111000010010101",
    "1111001110001101",
    "1111011101111101",
    "1111110000101011",
    "1111111010110111",
    "1111100110011101",
    "1111010100000110",
    "1111000101101010",
    "1110111100010100",
    "1110111000001110",
    "1110111000011101",
    "1110111011011000",
    "1110111111001100",
    "1111000010100111",
    "1111000100110110",
    "1111000101110001",
    "1111000101100010",
    "1111000100011100",
    "1111000010101011",
    "1111000000001101",
    "1110111101000100",
    "1110111001010000",
    "1110110100111011",
    "1110110000011111",
    "1110101100011100",
    "1110101001010101",
    "1110100111100011",
    "1110100111011010",
    "1110101001000010",
    "1110101100011110",
    "1110110001100110",
    "1110111000001100",
    "1110111111111000",
    "1111001000001000",
    "1111010000010101",
    "1111011000000110",
    "1111011110111111",
    "1111100101001000",
    "1111101011100000",
    "1111110011111111",
    "1111111111100001",
    "1111101101111011",
    "1111010111011010",
    "1110111101110000",
    "1110100011111100",
    "1110001101010001",
    "1101111100010011",
    "1101110010000011",
    "1101101110001111",
    "1101101111011001",
    "1101110011100110",
    "1101111001000001",
    "1101111110010111",
    "1110000010111001",
    "1110000110010101",
    "1110001000110000",
    "1110001010001110",
    "1110001010110000",
    "1110001010011001",
    "1110001001001100",
    "1110000111010101",
    "1110000101001000",
    "1110000011000000",
    "1110000001010101",
    "1110000000100001",
    "1110000000111001",
    "1110000010101111",
    "1110000110001000",
    "1110001010111100",
    "1110010001000010",
    "1110011000111010",
    "1110100100011101",
    "1110110101111110",
    "1111001110100110",
    "1111101101010100",
    "1111110001010101",
    "1111010010011100",
    "1110111010111101",
    "1110101110010100",
    "1110101100111100",
    "1110110100001101",
    "1111000000000000",
    "1111001100001010",
    "1111010101110110",
    "1111011100001110",
    "1111011111111111",
    "1111100010110011",
    "1111100110010011",
    "1111101010111101",
    "1111110000001111",
    "1111110100111100",
    "1111110111111000",
    "1111111000101011",
    "1111110111111001",
    "1111110110110010",
    "1111110110100001",
    "1111110111110101",
    "1111111010111100",
    "1111111111100110",
    "1111111010101010",
    "1111110100100011",
    "1111101110100101",
    "1111101001000100",
    "1111100100001101",
    "1111100000000010",
    "1111011100101000",
    "1111011010001001",
    "1111011000111001",
    "1111011001001100",
    "1111011011100000",
    "1111100000000011",
    "1111100110101110",
    "1111101110111000",
    "1111110111011011",
    "1111111111000000",
    "1111111011110000",
    "1111111001101101",
    "1111111010100010",
    "1111111100111011",
    "1111111111000000",
    "1111111111001001",
    "1111111100101110",
    "1111111000001001",
    "1111110010100011",
    "1111101101000111",
    "1111101000101000",
    "1111100101010010",
    "1111100010110001",
    "1111100000100111",
    "1111011110011100",
    "1111011100001010",
    "1111011001111001",
    "1111010111111001",
    "1111010110001011",
    "1111010100101001",
    "1111010010111011",
    "1111010000110000",
    "1111001101111101",
    "1111001010101010",
    "1111000111011000",
    "1111000101000000",
    "1111000100010101",
    "1111000101101110",
    "1111001000110111",
    "1111001100110011",
    "1111010000010101",
    "1111010010010100",
    "1111010010000110",
    "1111001111111101",
    "1111001100110011",
    "1111001001111010",
    "1111001000001011",
    "1111000111110111",
    "1111001000011010",
    "1111001000111111",
    "1111001000111001",
    "1111000111110101",
    "1111000110010101",
    "1111000101010000",
    "1111000101100101",
    "1111000111111111",
    "1111001100100011",
    "1111010010110011",
    "1111011001111001",
    "1111100000111011",
    "1111100111010000",
    "1111101100101001",
    "1111110001011001",
    "1111110110010100",
    "1111111100001001",
    "1111111100101100",
    "1111110100101110",
    "1111101101000011",
    "1111100111000100",
    "1111100011110100",
    "1111100011100001",
    "1111100101001110",
    "1111100111011100",
    "1111101000100010",
    "1111100111101000",
    "1111100100111011",
    "1111100001101001",
    "1111011111011001",
    "1111011111100100",
    "1111100010110100",
    "1111101001000011",
    "1111110001010100",
    "1111111010010101",
    "1111111101000111",
    "1111110101111101",
    "1111110000011111",
    "1111101100101001",
    "1111101010000111",
    "1111101000101101",
    "1111101000100011",
    "1111101001111111",
    "1111101101011011",
    "1111110010111001",
    "1111111001111100",
    "1111111110010000",
    "1111110110110101",
    "1111110000110110",
    "1111101101001000",
    "1111101100010011",
    "1111101110100000",
    "1111110011100000",
    "1111111010100111",
    "1111111101000110",
    "1111110100011110",
    "1111101011101111",
    "1111100010101100",
    "1111011001001100",
    "1111001111101001",
    "1111000111010000",
    "1111000001100110",
    "1111000000000111",
    "1111000011010010",
    "1111001010010011",
    "1111010011010010",
    "1111011100001110",
    "1111100011100010",
    "1111101000100010",
    "1111101011010110",
    "1111101100100101",
    "1111101100110101",
    "1111101100100111",
    "1111101100001101",
    "1111101011111011",
    "1111101100001110",
    "1111101101100100",
    "1111110000011001",
    "1111110100110111",
    "1111111010110111",
    "1111111110000110",
    "1111110110111001",
    "1111110000011011",
    "1111101011101100",
    "1111101001100010",
    "1111101010100001",
    "1111101110011110",
    "1111110100100001",
    "1111111011000010",
    "1111111111110100",
    "1111111101101100",
    "1111111111001101",
    "1111111100000010",
    "1111110101011000",
    "1111101110011000",
    "1111101000010111",
    "1111100100000101",
    "1111100001110100",
    "1111100001101110",
    "1111100011111000",
    "1111101000010101",
    "1111101110111101",
    "1111110111000111",
    "1111111111100111",
    "1111111001000100",
    "1111110100101001",
    "1111110100010000",
    "1111111000011000",
    "1111111111010000",
    "1111110011110010",
    "1111100110111101",
    "1111011010111100",
    "1111010001110100",
    "1111001101001110",
    "1111001101111101",
    "1111010011111000",
    "1111011101111111",
    "1111101010101000",
    "1111110111101111",
    "1111111100011111",
    "1111110011011001",
    "1111101101011011",
    "1111101010011001",
    "1111101001101100",
    "1111101010100100",
    "1111101100100100",
    "1111101111100110",
    "1111110011100111",
    "1111111000010111",
    "1111111100111111",
    "1111111111110000",
    "1111111111000101",
    "1111111110011110",
    "1111111001001111",
    "1111110010000111",
    "1111101010001111",
    "1111100010101011",
    "1111011100001100",
    "1111010111011000",
    "1111010100100000",
    "1111010011101111",
    "1111010100111110",
    "1111011000000011",
    "1111011100110101",
    "1111100011011000",
    "1111101011111010",
    "1111110110011110",
    "1111111101010110",
    "1111110000100110",
    "1111100100101001",
    "1111011010100011",
    "1111010010110110",
    "1111001101001111",
    "1111001001000001",
    "1111000101100000",
    "1111000010100001",
    "1111000000010001",
    "1110111111010111",
    "1111000000010001",
    "1111000011001101",
    "1111001000000011",
    "1111001110011011",
    "1111010101110111",
    "1111011101111011",
    "1111100110001000",
    "1111101101110111",
    "1111110100100011",
    "1111111001011101",
    "1111111011111100",
    "1111111011100001",
    "1111111000000001",
    "1111110001101011",
    "1111101001001010",
    "1111011111011100",
    "1111010101110010",
    "1111001101100011",
    "1111000111111100",
    "1111000110000001",
    "1111001000010011",
    "1111001110101000",
    "1111011000010000",
    "1111100011111100",
    "1111110000011100",
    "1111111100101010",
    "1111110111111110",
    "1111101101110010",
    "1111100100110011",
    "1111011100111111",
    "1111010110011111",
    "1111010001010100",
    "1111001101100011",
    "1111001010111010",
    "1111001000111100",
    "1111000111000100",
    "1111000100110001",
    "1111000001101110",
    "1110111101110101",
    "1110111001010101",
    "1110110100101111",
    "1110110000101110",
    "1110101101101110",
    "1110101100000100",
    "1110101011101010",
    "1110101100001110",
    "1110101101010100",
    "1110101110101000",
    "1110101111110110",
    "1110110001000000",
    "1110110010001000",
    "1110110011011000",
    "1110110100111011",
    "1110110110110110",
    "1110111001001100",
    "1110111100000010",
    "1110111111010100",
    "1111000010111110",
    "1111000110111011",
    "1111001011000111",
    "1111001111100001",
    "1111010100000110",
    "1111011000110000",
    "1111011101011011",
    "1111100001111110",
    "1111100110111010",
    "1111101101111011",
    "1111111001101111",
    "1111110011010011",
    "1111011000110000",
    "1110111000111100",
    "1110011000100011",
    "1101111101010010",
    "1101101011110101",
    "1101100110000100",
    "1101101010011011",
    "1101110100101111",
    "1110000000000010",
    "1110001000011110",
    "1110001100011100",
    "1110001100010110",
    "1110001001111100",
    "1110000111001101",
    "1110000101011111",
    "1110000101000110",
    "1110000101101001",
    "1110000110010011",
    "1110000110101000",
    "1110000110101000",
    "1110000110100111",
    "1110000110110100",
    "1110000111010101",
    "1110001000000110",
    "1110001001101111",
    "1110001110011011",
    "1110011001010101",
    "1110101100101000",
    "1111001000001011",
    "1111101000111000",
    "1111110110011100",
    "1111011011011011",
    "1111001010001111",
    "1111000100000110",
    "1111000110110001",
    "1111001110001010",
    "1111010110010110",
    "1111011100111100",
    "1111100001101011",
    "1111100101101111",
    "1111101010100010",
    "1111110000111000",
    "1111111000001110",
    "1111111111000100",
    "1111111100000001",
    "1111111001111001",
    "1111111010010010",
    "1111111100001010",
    "1111111110001110",
    "1111111111101101",
    "1111111111101100",
    "1111111111111000",
    "1111111110011110",
    "1111111011111001",
    "1111110111111111",
    "1111110010101010",
    "1111101100000000",
    "1111100100010111",
    "1111011100010011",
    "1111010100100100",
    "1111001101111000",
    "1111001000110010",
    "1111000101100101",
    "1111000100010111",
    "1111000100111110",
    "1111000111010101",
    "1111001011010001",
    "1111010000101001",
    "1111010111001011",
    "1111011110010110",
    "1111100101101001",
    "1111101100111001",
    "1111110100001010",
    "1111111011100100",
    "1111111101000001",
    "1111110110010011",
    "1111110001000010",
    "1111101101101110",
    "1111101100010111",
    "1111101100010001",
    "1111101100100010",
    "1111101100011011",
    "1111101011101011",
    "1111101010100011",
    "1111101001100110",
    "1111101001011001",
    "1111101010001111",
    "1111101011111101",
    "1111101101111100",
    "1111101111010111",
    "1111101111011010",
    "1111101101100100",
    "1111101001101010",
    "1111100100001011",
    "1111011101111101",
    "1111010111111111",
    "1111010010111101",
    "1111001110111111",
    "1111001011110011",
    "1111001000110010",
    "1111000101011011",
    "1111000001101100",
    "1110111110000100",
    "1110111011010100",
    "1110111010000111",
    "1110111010101101",
    "1110111100101011",
    "1110111111010001",
    "1111000001101110",
    "1111000011101111",
    "1111000101011111",
    "1111000111100010",
    "1111001010011101",
    "1111001110010110",
    "1111010010101110",
    "1111010110101111",
    "1111011001101111",
    "1111011011100000",
    "1111011100100001",
    "1111011101101101",
    "1111100000000111",
    "1111100100011100",
    "1111101010110000",
    "1111110010010011",
    "1111111001110010",
    "1111111111101101",
    "1111111101001111",
    "1111111101110001",
    "1111111110011110",
    "1111111001000001",
    "1111110100000000",
    "1111110001100111",
    "1111110011000111",
    "1111111000011001",
    "1111111111111010",
    "1111110111111111",
    "1111110001110010",
    "1111101110100011",
    "1111101110100101",
    "1111110001010100",
    "1111110101110100",
    "1111111011001011",
    "1111111111001001",
    "1111111001011110",
    "1111110011110010",
    "1111101110001110",
    "1111101001001111",
    "1111100101100010",
    "1111100011110011",
    "1111100100011101",
    "1111100111010110",
    "1111101011101110",
    "1111110000100100",
    "1111110100111001",
    "1111110111110110",
    "1111111000111000",
    "1111110111101000",
    "1111110100000111",
    "1111101110110001",
    "1111101000011110",
    "1111100010010100",
    "1111011101001100",
    "1111011001011011",
    "1111010110101111",
    "1111010100100010",
    "1111010010010010",
    "1111001111101110",
    "1111001100111000",
    "1111001010000001",
    "1111000111010011",
    "1111000100111001",
    "1111000010111001",
    "1111000001100110",
    "1111000001010111",
    "1111000010101011",
    "1111000101110100",
    "1111001010111010",
    "1111010001110001",
    "1111011001111010",
    "1111100010100100",
    "1111101010101011",
    "1111110001000010",
    "1111110100101010",
    "1111110100111111",
    "1111110010010000",
    "1111101101100010",
    "1111101000100000",
    "1111100101000001",
    "1111100100101001",
    "1111101000001001",
    "1111101111100010",
    "1111111010000111",
    "1111111001000101",
    "1111101011010011",
    "1111011101101001",
    "1111010001001010",
    "1111000110110110",
    "1110111111101100",
    "1110111100100110",
    "1110111101111111",
    "1111000011101110",
    "1111001100111100",
    "1111011000010000",
    "1111100100000101",
    "1111101111000000",
    "1111111000000110",
    "1111111110111011",
    "1111111100011110",
    "1111111001111111",
    "1111111001011110",
    "1111111010110011",
    "1111111101110111",
    "1111111101100001",
    "1111110111110011",
    "1111110001010101",
    "1111101010101001",
    "1111100100001101",
    "1111011110100001",
    "1111011001111111",
    "1111010110111001",
    "1111010101010000",
    "1111010100111011",
    "1111010101011111",
    "1111010110011011",
    "1111010111010001",
    "1111010111111010",
    "1111011000100101",
    "1111011001110100",
    "1111011100010001",
    "1111100000010010",
    "1111100101110100",
    "1111101100100100",
    "1111110100000011",
    "1111111011110110",
    "1111111100010111",
    "1111110100111000",
    "1111101110000011",
    "1111101000011001",
    "1111100100010111",
    "1111100010000000",
    "1111100001000011",
    "1111100000110110",
    "1111100000111001",
    "1111100001000010",
    "1111100001010100",
    "1111100001110110",
    "1111100010011111",
    "1111100010110110",
    "1111100010101001",
    "1111100001111011",
    "1111100001011010",
    "1111100010010101",
    "1111100110000011",
    "1111101101011010",
    "1111111000011011",
    "1111111001110000",
    "1111101010110010",
    "1111011100011100",
    "1111010000011110",
    "1111001000000011",
    "1111000011111000",
    "1111000100000000",
    "1111000111111001",
    "1111001110011110",
    "1111010110010101",
    "1111011110000000",
    "1111100100001011",
    "1111101000000000",
    "1111101001001100",
    "1111100111110110",
    "1111100100010010",
    "1111011110111011",
    "1111011000010000",
    "1111010000111001",
    "1111001001101111",
    "1111000011110100",
    "1111000000001100",
    "1110111111101001",
    "1111000010101011",
    "1111001001000010",
    "1111010010010100",
    "1111011101101011",
    "1111101010010000",
    "1111110111000111",
    "1111111100101110",
    "1111110010010110",
    "1111101010100001",
    "1111100101101110",
    "1111100011111100",
    "1111100100101100",
    "1111100111000011",
    "1111101001111110",
    "1111101100100110",
    "1111101110010000",
    "1111101110101001",
    "1111101101101111",
    "1111101011100110",
    "1111101000010011",
    "1111100100000110",
    "1111011111001101",
    "1111011001111010",
    "1111010100010101",
    "1111001110101101",
    "1111001001000110",
    "1111000011101110",
    "1110111110110110",
    "1110111010101111",
    "1110110111100011",
    "1110110101011111",
    "1110110100100100",
    "1110110100101001",
    "1110110101011101",
    "1110110110101100",
    "1110111000000011",
    "1110111001010011",
    "1110111010100000",
    "1110111011110000",
    "1110111101010010",
    "1110111111010100",
    "1111000001111000",
    "1111000100110110",
    "1111001000000001",
    "1111001011001111",
    "1111001110011100",
    "1111010001101011",
    "1111010100111110",
    "1111011000011110",
    "1111011100001010",
    "1111100000000010",
    "1111100100000000",
    "1111101000000111",
    "1111101101000000",
    "1111110100101101",
    "1111111101111110",
    "1111101000111110",
    "1111001100001110",
    "1110101010100110",
    "1110001001010000",
    "1101101101111010",
    "1101011101000100",
    "1101011000010000",
    "1101011101100001",
    "1101101000100111",
    "1101110100100111",
    "1101111101110111",
    "1110000010110011",
    "1110000011110001",
    "1110000010010100",
    "1110000000010001",
    "1101111110101110",
    "1101111110000010",
    "1101111101111000",
    "1101111101110000",
    "1101111101011110",
    "1101111101010010",
    "1101111101101011",
    "1101111110111010",
    "1110000000111000",
    "1110000011010011",
    "1110000110000001",
    "1110001001000111",
    "1110001101001110",
    "1110010100000101",
    "1110100000001000",
    "1110110011000110",
    "1111001100110010",
    "1111101010100110",
    "1111110111100101",
    "1111011110010110",
    "1111001101001111",
    "1111000101111011",
    "1111000111100111",
    "1111001111110001",
    "1111011011010011",
    "1111100111010101",
    "1111110001110010",
    "1111111001010111",
    "1111111101100011",
    "1111111110100100",
    "1111111101001000",
    "1111111010001010",
    "1111110110100111",
    "1111110011010101",
    "1111110001001000",
    "1111110000110001",
    "1111110010111101",
    "1111110111110101",
    "1111111110111011",
    "1111111000101101",
    "1111110000001111",
    "1111101000101011",
    "1111100010111011",
    "1111011111101011",
    "1111011111001000",
    "1111100001000000",
    "1111100100010111",
    "1111101000000011",
    "1111101010111101",
    "1111101100001101",
    "1111101011011110",
    "1111101000111011",
    "1111100101011000",
    "1111100010000011",
    "1111100000010101",
    "1111100001011010",
    "1111100101101110",
    "1111101100101011",
    "1111110100110110",
    "1111111100100001",
    "1111111101011101",
    "1111111001011000",
    "1111110110100001",
    "1111110011110110",
    "1111110000100011",
    "1111101100010011",
    "1111100111010000",
    "1111100001110011",
    "1111011100010110",
    "1111010111001101",
    "1111010010101111",
    "1111001111010001",
    "1111001101000100",
    "1111001100010001",
    "1111001100101010",
    "1111001101101000",
    "1111001110010111",
    "1111001110001010",
    "1111001100100101",
    "1111001001101111",
    "1111000110000011",
    "1111000010001010",
    "1110111110110001",
    "1110111100010100",
    "1110111010111111",
    "1110111010100101",
    "1110111010110101",
    "1110111011010100",
    "1110111011100001",
    "1110111011001100",
    "1110111010001111",
    "1110111000111100",
    "1110110111110010",
    "1110110111010101",
    "1110111000001001",
    "1110111010011000",
    "1110111101111000",
    "1111000010010010",
    "1111000111000110",
    "1111001011110011",
    "1111010000001100",
    "1111010100000011",
    "1111010111010101",
    "1111011001111111",
    "1111011100000101",
    "1111011101110011",
    "1111011111010100",
    "1111100001000010",
    "1111100011010010",
    "1111100110010101",
    "1111101010001111",
    "1111101110110011",
    "1111110011110010",
    "1111111000111111",
    "1111111110010010",
    "1111111100001111",
    "1111110110110011",
    "1111110001101010",
    "1111101101011000",
    "1111101010100011",
    "1111101001101001",
    "1111101010110010",
    "1111101101101011",
    "1111110001101100",
    "1111110110001010",
    "1111111010100011",
    "1111111110110101",
    "1111111100110010",
    "1111111000001001",
    "1111110011001111",
    "1111101110010010",
    "1111101001101101",
    "1111100110001000",
    "1111100100001000",
    "1111100100001101",
    "1111100110110101",
    "1111101100010101",
    "1111110100100100",
    "1111111110110111",
    "1111110110001000",
    "1111101100001100",
    "1111100100110110",
    "1111100001001111",
    "1111100001101001",
    "1111100101110100",
    "1111101101001110",
    "1111110111010011",
    "1111111100001111",
    "1111101101111000",
    "1111011110010110",
    "1111001110111000",
    "1111000001000111",
    "1110110110100101",
    "1110110000100001",
    "1110101111011010",
    "1110110011000011",
    "1110111010100010",
    "1111000100101010",
    "1111001111111101",
    "1111011010111100",
    "1111100100010101",
    "1111101011001111",
    "1111101111001001",
    "1111101111111101",
    "1111101101111001",
    "1111101001100000",
    "1111100011101001",
    "1111011101010110",
    "1111010111111010",
    "1111010100101100",
    "1111010100111011",
    "1111011001010011",
    "1111100001111000",
    "1111101101110111",
    "1111111011110110",
    "1111110101111010",
    "1111101001010011",
    "1111011111110001",
    "1111011010011011",
    "1111011001101011",
    "1111011101011100",
    "1111100100110011",
    "1111101110010110",
    "1111111000001111",
    "1111111111011001",
    "1111111010000111",
    "1111111000101000",
    "1111111010101101",
    "1111111111010101",
    "1111111010101101",
    "1111110100100000",
    "1111101110101001",
    "1111101001011101",
    "1111100101010010",
    "1111100010101110",
    "1111100010011111",
    "1111100101000001",
    "1111101010010000",
    "1111110001010100",
    "1111111000110001",
    "1111111111000101",
    "1111111101000001",
    "1111111100010001",
    "1111111110100111",
    "1111111100011110",
    "1111110110000001",
    "1111101111000111",
    "1111101001000001",
    "1111100100101110",
    "1111100010111101",
    "1111100011111100",
    "1111100111011110",
    "1111101100110000",
    "1111110010110010",
    "1111111000100010",
    "1111111101010100",
    "1111111111000101",
    "1111111100011111",
    "1111111010011001",
    "1111111000011001",
    "1111110110001111",
    "1111110011111000",
    "1111110001010011",
    "1111101110011010",
    "1111101011001010",
    "1111100111101001",
    "1111100100001010",
    "1111100001001000",
    "1111011110111011",
    "1111011101101011",
    "1111011101001001",
    "1111011100111111",
    "1111011100111101",
    "1111011101001110",
    "1111011110010100",
    "1111100000111101",
    "1111100101110110",
    "1111101101010001",
    "1111110110111110",
    "1111111101110001",
    "1111110010010011",
    "1111100111111110",
    "1111011111111010",
    "1111011010101101",
    "1111011000010110",
    "1111011000000011",
    "1111011000101000",
    "1111011000110111",
    "1111010111101100",
    "1111010100101010",
    "1111010000000011",
    "1111001010100101",
    "1111000101010000",
    "1111000000111011",
    "1110111101111011",
    "1110111100001100",
    "1110111011001111",
    "1110111010110100",
    "1110111010110111",
    "1110111100000101",
    "1110111111011111",
    "1111000110000110",
    "1111010000010100",
    "1111011101100011",
    "1111101100001101",
    "1111111010000100",
    "1111111010111110",
    "1111110100011001",
    "1111110010100101",
    "1111110100111110",
    "1111111010011000",
    "1111111110100010",
    "1111110111001000",
    "1111110000011110",
    "1111101011011101",
    "1111101000101100",
    "1111101000100001",
    "1111101011000000",
    "1111101111111100",
    "1111110111000011",
    "1111111111110100",
    "1111110110010101",
    "1111101100010100",
    "1111100010111001",
    "1111011010110100",
    "1111010100010101",
    "1111001111011010",
    "1111001011101010",
    "1111001000101010",
    "1111000110001011",
    "1111000100010011",
    "1111000011011000",
    "1111000011101110",
    "1111000101010101",
    "1111000111110001",
    "1111001010001001",
    "1111001011011101",
    "1111001011000010",
    "1111001000110101",
    "1111000101100010",
    "1111000010001101",
    "1110111111111010",
    "1110111111000111",
    "1110111111110011",
    "1111000001010100",
    "1111000010111011",
    "1111000100001011",
    "1111000101000000",
    "1111000101110100",
    "1111000111001001",
    "1111001001100011",
    "1111001101001111",
    "1111010010000110",
    "1111010111101101",
    "1111011101100001",
    "1111100011000011",
    "1111100111111011",
    "1111101100000101",
    "1111101111110001",
    "1111110100101100",
    "1111111110001101",
    "1111110000011110",
    "1111010110011000",
    "1110110101101110",
    "1110010011101111",
    "1101110110110100",
    "1101100100011100",
    "1101011111000111",
    "1101100101001001",
    "1101110001101011",
    "1101111110110110",
    "1110001000001100",
    "1110001011110111",
    "1110001010011101",
    "1110000110000001",
    "1110000000111110",
    "1101111101000100",
    "1101111010101000",
    "1101111001011000",
    "1101111000101010",
    "1101111000000110",
    "1101111000000100",
    "1101111001001110",
    "1101111011111100",
    "1101111111111101",
    "1110000100101001",
    "1110001001100010",
    "1110001111001100",
    "1110010111010001",
    "1110100011100010",
    "1110110100111100",
    "1111001010111010",
    "1111100011001101",
    "1111111010101010",
    "1111110001111001",
    "1111100100101110",
    "1111011110000101",
    "1111011100110101",
    "1111011110110110",
    "1111100010010000",
    "1111100101111100",
    "1111101001100011",
    "1111101101001001",
    "1111110000110010",
    "1111110100001001",
    "1111110110100110",
    "1111110111110000",
    "1111110111110100",
    "1111110111100010",
    "1111110111111001",
    "1111111001100101",
    "1111111100101010",
    "1111111111010111",
    "1111111011010011",
    "1111110111101100",
    "1111110100100101",
    "1111110001100111",
    "1111101110010001",
    "1111101010001001",
    "1111100101010000",
    "1111100000000010",
    "1111011010111100",
    "1111010110010000",
    "1111010010000110",
    "1111001110011100",
    "1111001011011011",
    "1111001001100101",
    "1111001001101010",
    "1111001100011110",
    "1111010010100001",
    "1111011011100001",
    "1111100110100100",
    "1111110010010110",
    "1111111101101010",
    "1111111000010001",
    "1111101111110110",
    "1111101001000011",
    "1111100011110100",
    "1111100000000101",
    "1111011101111010",
    "1111011101010010",
    "1111011110001001",
    "1111100000011001",
    "1111100011110001",
    "1111101000000111",
    "1111101100111010",
    "1111110001011111",
    "1111110101000011",
    "1111110110110010",
    "1111110110010101",
    "1111110011101100",
    "1111101111010100",
    "1111101001111010",
    "1111100100000101",
    "1111011110000010",
    "1111010111101100",
    "1111010000110001",
    "1111001001001100",
    "1111000001010100",
    "1110111001110111",
    "1110110011110110",
    "1110110000000111",
    "1110101111001100",
    "1110110000111101",
    "1110110100110100",
    "1110111001111100",
    "1110111111010100",
    "1111000100000000",
    "1111000111010000",
    "1111001000100011",
    "1111000111110010",
    "1111000101010010",
    "1111000001111101",
    "1110111110111101",
    "1110111101011100",
    "1110111110001101",
    "1111000001011110",
    "1111000110110100",
    "1111001101100100",
    "1111010100110100",
    "1111011011101111",
    "1111100001100111",
    "1111100110000011",
    "1111101000110101",
    "1111101010000111",
    "1111101010010101",
    "1111101001111101",
    "1111101001100000",
    "1111101001011011",
    "1111101010000010",
    "1111101011101110",
    "1111101110111000",
    "1111110011110001",
    "1111111010011001",
    "1111111101110011",
    "1111110110000001",
    "1111101111101011",
    "1111101100001010",
    "1111101100011011",
    "1111110000110000",
    "1111111000100111",
    "1111111101000111",
    "1111110001111111",
    "1111100111100000",
    "1111011110110110",
    "1111011001000010",
    "1111010110100111",
    "1111010111110010",
    "1111011100010111",
    "1111100011101111",
    "1111101100110111",
    "1111110110011000",
    "1111111110110010",
    "1111111011001100",
    "1111111000100100",
    "1111111001101111",
    "1111111110100100",
    "1111111001011100",
    "1111101111010111",
    "1111100100011111",
    "1111011010010001",
    "1111010001111001",
    "1111001100001001",
    "1111001001001001",
    "1111001000010110",
    "1111001000111001",
    "1111001001111010",
    "1111001010111010",
    "1111001011110010",
    "1111001100100110",
    "1111001101011110",
    "1111001110001111",
    "1111001110100100",
    "1111001110001010",
    "1111001100110011",
    "1111001010101101",
    "1111001000010110",
    "1111000110011011",
    "1111000101101010",
    "1111000110100111",
    "1111001001100010",
    "1111001110010010",
    "1111010100100100",
    "1111011011101101",
    "1111100011000000",
    "1111101001110001",
    "1111101111011100",
    "1111110011110110",
    "1111110110111111",
    "1111111001001100",
    "1111111010111001",
    "1111111100101010",
    "1111111111000000",
    "1111111101100110",
    "1111111000111101",
    "1111110011000001",
    "1111101100000000",
    "1111100100010101",
    "1111011100101101",
    "1111010110001000",
    "1111010001101011",
    "1111010000010010",
    "1111010010010100",
    "1111010111010101",
    "1111011110001010",
    "1111100101011000",
    "1111101011110110",
    "1111110001000110",
    "1111110101010111",
    "1111111001001010",
    "1111111100111011",
    "1111111111011011",
    "1111111100100001",
    "1111111011010010",
    "1111111100011100",
    "1111111111100110",
    "1111111001001011",
    "1111110000111001",
    "1111100111110001",
    "1111011110110110",
    "1111010111001101",
    "1111010001100001",
    "1111001110001010",
    "1111001100111111",
    "1111001101011110",
    "1111001110110101",
    "1111010000010101",
    "1111010001101001",
    "1111010010111101",
    "1111010101000001",
    "1111011000111010",
    "1111011111010110",
    "1111101000010110",
    "1111110011001010",
    "1111111110011111",
    "1111110111000100",
    "1111101110100011",
    "1111101000011100",
    "1111100100101001",
    "1111100010101111",
    "1111100010001101",
    "1111100010011100",
    "1111100011000001",
    "1111100011100010",
    "1111100011110001",
    "1111100011101111",
    "1111100011110001",
    "1111100100001010",
    "1111100101010011",
    "1111100111011010",
    "1111101010011100",
    "1111101110001101",
    "1111110010010101",
    "1111110110010101",
    "1111111001110001",
    "1111111100011010",
    "1111111110011001",
    "1111111111100110",
    "1111111100110001",
    "1111111000001011",
    "1111110001010111",
    "1111101000100011",
    "1111011110101000",
    "1111010100111011",
    "1111001100101101",
    "1111000110110001",
    "1111000011000110",
    "1111000001000101",
    "1110111111101001",
    "1110111101111111",
    "1110111011101011",
    "1110111001001011",
    "1110110111011000",
    "1110110111100101",
    "1110111010110101",
    "1111000001100110",
    "1111001011100110",
    "1111010111111001",
    "1111100100111110",
    "1111110001001100",
    "1111111011001010",
    "1111111110000010",
    "1111111010101010",
    "1111111010001101",
    "1111111011101000",
    "1111111101110001",
    "1111111111100010",
    "1111111111110001",
    "1111111111100000",
    "1111111101101001",
    "1111111011000001",
    "1111111000001000",
    "1111110101011000",
    "1111110010111111",
    "1111110001000010",
    "1111101111011110",
    "1111101110001000",
    "1111101100110111",
    "1111101011100011",
    "1111101010000010",
    "1111101000010100",
    "1111100110011110",
    "1111100100101001",
    "1111100011000101",
    "1111100010000010",
    "1111100001101001",
    "1111100001110011",
    "1111100010000010",
    "1111100001101110",
    "1111100000001101",
    "1111011101001010",
    "1111011000100011",
    "1111010010110110",
    "1111001100110101",
    "1111000111011011",
    "1111000011011010",
    "1111000001001111",
    "1111000000110110",
    "1111000001111011",
    "1111000011110110",
    "1111000110000110",
    "1111001000010001",
    "1111001010010011",
    "1111001100010111",
    "1111001110101101",
    "1111010001100110",
    "1111010101000101",
    "1111011001000010",
    "1111011101010010",
    "1111100001100001",
    "1111100101100000",
    "1111101001001100",
    "1111101100101010",
    "1111110000100001",
    "1111110110100110",
    "1111111110010010",
    "1111101011111010",
    "1111010001101110",
    "1110110010000101",
    "1110010001100110",
    "1101110101101110",
    "1101100011000011",
    "1101011011100011",
    "1101011101110011",
    "1101100101111100",
    "1101101111010100",
    "1101110110010000",
    "1101111001010000",
    "1101111000101010",
    "1101110110001101",
    "1101110011111000",
    "1101110011000011",
    "1101110100001101",
    "1101110110111100",
    "1101111010100101",
    "1101111110010111",
    "1110000010000011",
    "1110000101100010",
    "1110001000101101",
    "1110001011001111",
    "1110001100111101",
    "1110001101110101",
    "1110001110010111",
    "1110001111010100",
    "1110010001111011",
    "1110011000010110",
    "1110100100111001",
    "1110111000101100",
    "1111010010110001",
    "1111101111111011",
    "1111110100010110",
    "1111011110101101",
    "1111010010010101",
    "1111010000000010",
    "1111010101111001",
    "1111100000010001",
    "1111101011001110",
    "1111110011110111",
    "1111111000110011",
    "1111111010001001",
    "1111111001000001",
    "1111110111000000",
    "1111110101011110",
    "1111110101000110",
    "1111110101110111",
    "1111110111011000",
    "1111111001010110",
    "1111111011110001",
    "1111111110111000",
    "1111111101010001",
    "1111111001000101",
    "1111110101000111",
    "1111110001111101",
    "1111110000000001",
    "1111101111100000",
    "1111110000010111",
    "1111110010001001",
    "1111110100001010",
    "1111110101100100",
    "1111110101101110",
    "1111110100010010",
    "1111110001001101",
    "1111101100111011",
    "1111101000010011",
    "1111100100101001",
    "1111100011011000",
    "1111100101101110",
    "1111101100000111",
    "1111110110010000",
    "1111111101001001",
    "1111110000000000",
    "1111100100001000",
    "1111011010111000",
    "1111010100111011",
    "1111010010010100",
    "1111010010110110",
    "1111010110000100",
    "1111011011001100",
    "1111100000111101",
    "1111100101110010",
    "1111101000001111",
    "1111100111010010",
    "1111100010110001",
    "1111011011011011",
    "1111010010101001",
    "1111001010001110",
    "1111000011101001",
    "1110111111110011",
    "1110111110101101",
    "1110111111100100",
    "1111000001000111",
    "1111000001111001",
    "1111000000110110",
    "1110111101100001",
    "1110111000010110",
    "1110110010011010",
    "1110101101000100",
    "1110101001100010",
    "1110101000100010",
    "1110101010001001",
    "1110101101110011",
    "1110110010100100",
    "1110110111011101",
    "1110111011110101",
    "1110111111100011",
    "1111000010111000",
    "1111000110001000",
    "1111001001011110",
    "1111001100101000",
    "1111001110111101",
    "1111001111101011",
    "1111001110010111",
    "1111001011001001",
    "1111000110110010",
    "1111000010011111",
    "1110111111100001",
    "1110111111000010",
    "1111000001111000",
    "1111001000010110",
    "1111010010001111",
    "1111011110101000",
    "1111101100000101",
    "1111111000111001",
    "1111111100011101",
    "1111110101000110",
    "1111110001010011",
    "1111110000100111",
    "1111110010001100",
    "1111110101001001",
    "1111111000111101",
    "1111111101011010",
    "1111111101100011",
    "1111111000000110",
    "1111110010100110",
    "1111101101101000",
    "1111101001110101",
    "1111100111101000",
    "1111100111001001",
    "1111101000001111",
    "1111101010101110",
    "1111101110100010",
    "1111110011101110",
    "1111111010001001",
    "1111111110100010",
    "1111110111001100",
    "1111110000110000",
    "1111101100000111",
    "1111101001101101",
    "1111101001100001",
    "1111101011000100",
    "1111101101100111",
    "1111110000011001",
    "1111110010110100",
    "1111110100101010",
    "1111110110001010",
    "1111110111111101",
    "1111111011000101",
    "1111111111010011",
    "1111110110011111",
    "1111101010100011",
    "1111011100101000",
    "1111001110101011",
    "1111000010111001",
    "1110111010111010",
    "1110110111011011",
    "1110111000000100",
    "1110111011110010",
    "1111000001001000",
    "1111000111000001",
    "1111001100101110",
    "1111010010000101",
    "1111010111000011",
    "1111011011100110",
    "1111011111101000",
    "1111100010110100",
    "1111100100111011",
    "1111100101110010",
    "1111100101101010",
    "1111100101000000",
    "1111100100101001",
    "1111100101010101",
    "1111100111101100",
    "1111101011111100",
    "1111110001110101",
    "1111111000110001",
    "1111111111111000",
    "1111111001101011",
    "1111110100101111",
    "1111110001101010",
    "1111110000100001",
    "1111110001000101",
    "1111110011000000",
    "1111110101110010",
    "1111111000110011",
    "1111111011010110",
    "1111111100101011",
    "1111111100001001",
    "1111111001011101",
    "1111110100111010",
    "1111101111011101",
    "1111101010100000",
    "1111100111011100",
    "1111100111010000",
    "1111101010001011",
    "1111101111101010",
    "1111110110011011",
    "1111111100111011",
    "1111111110001100",
    "1111111011110111",
    "1111111100001101",
    "1111111110110100",
    "1111111100111101",
    "1111110111111001",
    "1111110010011111",
    "1111101100111010",
    "1111100111001001",
    "1111100001001000",
    "1111011010111100",
    "1111010100111100",
    "1111001111110011",
    "1111001100011001",
    "1111001011101101",
    "1111001110100001",
    "1111010101001011",
    "1111011111001111",
    "1111101011100100",
    "1111111000011011",
    "1111111011110010",
    "1111110010011001",
    "1111101011110111",
    "1111101000000111",
    "1111100110100110",
    "1111100110101011",
    "1111100111110101",
    "1111101001101000",
    "1111101011101010",
    "1111101101100010",
    "1111101110110100",
    "1111101111010110",
    "1111101111001000",
    "1111101110010111",
    "1111101101001110",
    "1111101011101110",
    "1111101001110101",
    "1111100111100111",
    "1111100101010011",
    "1111100011011000",
    "1111100010100110",
    "1111100011101001",
    "1111100111001101",
    "1111101101101110",
    "1111110111011010",
    "1111111011110010",
    "1111101100100011",
    "1111011100000010",
    "1111001011110011",
    "1110111101100110",
    "1110110010111000",
    "1110101100011100",
    "1110101010000111",
    "1110101010111010",
    "1110101101010110",
    "1110110000001010",
    "1110110010100110",
    "1110110100101111",
    "1110110111010101",
    "1110111011010110",
    "1111000001100111",
    "1111001010010110",
    "1111010101000000",
    "1111100000011111",
    "1111101011011100",
    "1111110100100000",
    "1111111010101000",
    "1111111101010010",
    "1111111100101000",
    "1111111001011010",
    "1111110100110111",
    "1111110000010000",
    "1111101100100011",
    "1111101010001000",
    "1111101000110010",
    "1111100111111111",
    "1111100111010101",
    "1111100110110010",
    "1111100110110001",
    "1111100111111100",
    "1111101010110111",
    "1111101111110101",
    "1111110110101010",
    "1111111110101101",
    "1111111000110111",
    "1111110001001001",
    "1111101010111010",
    "1111100110110011",
    "1111100101000011",
    "1111100101100000",
    "1111100111101000",
    "1111101010100000",
    "1111101101000101",
    "1111101110010010",
    "1111101101011001",
    "1111101010000111",
    "1111100100101110",
    "1111011101110010",
    "1111010110000011",
    "1111001110000111",
    "1111000110100000",
    "1110111111011110",
    "1110111001010110",
    "1110110100011100",
    "1110110001000011",
    "1110101111011100",
    "1110101111101001",
    "1110110001100001",
    "1110110100101100",
    "1110111000101101",
    "1110111101001010",
    "1111000001110110",
    "1111000110101010",
    "1111001011100001",
    "1111010000011001",
    "1111010101000011",
    "1111011001001011",
    "1111011100100011",
    "1111011111000111",
    "1111100000111001",
    "1111100010010000",
    "1111100011100010",
    "1111100101010010",
    "1111101001010000",
    "1111110010101100",
    "1111111011100101",
    "1111100000111011",
    "1110111111101110",
    "1110011101000100",
    "1101111111000101",
    "1101101010111100",
    "1101100011001010",
    "1101100110001101",
    "1101101111110000",
    "1101111010101111",
    "1110000011001000",
    "1110000111010110",
    "1110000111111010",
    "1110000110011000",
    "1110000100101111",
    "1110000100001011",
    "1110000100110110",
    "1110000110000110",
    "1110000111010000",
    "1110000111110101",
    "1110001000001011",
    "1110001000110010",
    "1110001010000110",
    "1110001011111111",
    "1110001110000101",
    "1110010000000101",
    "1110010010001111",
    "1110010101100111",
    "1110011011111101",
    "1110100111000011",
    "1110110111100101",
    "1111001100110101",
    "1111100100011000",
    "1111111010111111",
    "1111110010011111",
    "1111100110000011",
    "1111011111110000",
    "1111011110001111",
    "1111011111011100",
    "1111100001110001",
    "1111100100100100",
    "1111101000000100",
    "1111101100101100",
    "1111110010011010",
    "1111111000010010",
    "1111111100111000",
    "1111111110110010",
    "1111111101010111",
    "1111111000111100",
    "1111110010111010",
    "1111101101010001",
    "1111101001111111",
    "1111101010011111",
    "1111101111010010",
    "1111110111111111",
    "1111111100100000",
    "1111101111111100",
    "1111100100000101",
    "1111011010100101",
    "1111010100100000",
    "1111010010000110",
    "1111010010100100",
    "1111010100100100",
    "1111010110101111",
    "1111011000010000",
    "1111011001001001",
    "1111011010001110",
    "1111011100110011",
    "1111100010001000",
    "1111101010101011",
    "1111110101111110",
    "1111111101010000",
    "1111110000101101",
    "1111100101110111",
    "1111011101110011",
    "1111011000110100",
    "1111010110110100",
    "1111010111011101",
    "1111011010010011",
    "1111011110111101",
    "1111100101000000",
    "1111101011111100",
    "1111110010111111",
    "1111111001001000",
    "1111111101010110",
    "1111111110110001",
    "1111111100111101",
    "1111111000000001",
    "1111110000101011",
    "1111100111111011",
    "1111011110101101",
    "1111010101011111",
    "1111001100010011",
    "1111000010111001",
    "1110111001010011",
    "1110110000000000",
    "1110101000001110",
    "1110100011011111",
    "1110100011010000",
    "1110101000001000",
    "1110110001100010",
    "1110111101101101",
    "1111001010000001",
    "1111010011111001",
    "1111011001100011",
    "1111011010011000",
    "1111010110110110",
    "1111010000001000",
    "1111000111101111",
    "1110111110110011",
    "1110110110001000",
    "1110101110010001",
    "1110100111110100",
    "1110100011011000",
    "1110100001110110",
    "1110100100000001",
    "1110101010011101",
    "1110110101000011",
    "1111000011000001",
    "1111010010110001",
    "1111100010001010",
    "1111101110111111",
    "1111110111100100",
    "1111111010111111",
    "1111111001011000",
    "1111110011110010",
    "1111101011111010",
    "1111100011101100",
    "1111011100111100",
    "1111011001000001",
    "1111011000101101",
    "1111011100001100",
    "1111100010111110",
    "1111101100001011",
    "1111110110011110",
    "1111111111100001",
    "1111110111011000",
    "1111110010010101",
    "1111110001001001",
    "1111110011110111",
    "1111111001101101",
    "1111111110101100",
    "1111110111000101",
    "1111110000110111",
    "1111101100111001",
    "1111101011010101",
    "1111101011110110",
    "1111101101110101",
    "1111110000110001",
    "1111110100010110",
    "1111111000010010",
    "1111111100010011",
    "1111111111111100",
    "1111111101010100",
    "1111111100001001",
    "1111111101000000",
    "1111111111101010",
    "1111111001110100",
    "1111110001100111",
    "1111100111101110",
    "1111011101001111",
    "1111010011100100",
    "1111001011111111",
    "1111000111010001",
    "1111000101011111",
    "1111000101111110",
    "1111000111100111",
    "1111001001011001",
    "1111001010110100",
    "1111001011111000",
    "1111001101000101",
    "1111001111000000",
    "1111010001111101",
    "1111010101111001",
    "1111011010010110",
    "1111011110100011",
    "1111100001110011",
    "1111100011101001",
    "1111100011111011",
    "1111100010111110",
    "1111100001010100",
    "1111011111100110",
    "1111011110101000",
    "1111011110111101",
    "1111100000111110",
    "1111100100101001",
    "1111101001100111",
    "1111101111010101",
    "1111110101010101",
    "1111111011010110",
    "1111111110101000",
    "1111111000100110",
    "1111110010011101",
    "1111101100001111",
    "1111100110001000",
    "1111100000011001",
    "1111011011001100",
    "1111010110110001",
    "1111010011010011",
    "1111010001010010",
    "1111010001010111",
    "1111010100001010",
    "1111011001111100",
    "1111100010011010",
    "1111101100101001",
    "1111110111001100",
    "1111111111011111",
    "1111111000110100",
    "1111110101100100",
    "1111110101111100",
    "1111111001101011",
    "1111111111101100",
    "1111110110111010",
    "1111101100100000",
    "1111100001000111",
    "1111010101011000",
    "1111001010000111",
    "1111000000001101",
    "1110111000100101",
    "1110110011111100",
    "1110110010101011",
    "1110110100110100",
    "1110111010000111",
    "1111000010001101",
    "1111001100100011",
    "1111011000100101",
    "1111100101011111",
    "1111110010001001",
    "1111111101010011",
    "1111111010001110",
    "1111110101010000",
    "1111110011110101",
    "1111110101010111",
    "1111111000101000",
    "1111111100010100",
    "1111111111001100",
    "1111111111100000",
    "1111111111110011",
    "1111111101010110",
    "1111111001011110",
    "1111110100101100",
    "1111101111011110",
    "1111101010000011",
    "1111100100100100",
    "1111011111001100",
    "1111011010001100",
    "1111010110000001",
    "1111010011010000",
    "1111010010100001",
    "1111010100010111",
    "1111011001000110",
    "1111100000110110",
    "1111101011010110",
    "1111110111111101",
    "1111111010011010",
    "1111101101010000",
    "1111100001111101",
    "1111011001100011",
    "1111010100011111",
    "1111010010010111",
    "1111010010001010",
    "1111010010100001",
    "1111010010010010",
    "1111010000101100",
    "1111001101110101",
    "1111001010010001",
    "1111000111000001",
    "1111000100111100",
    "1111000100101110",
    "1111000110011011",
    "1111001001111010",
    "1111001110100110",
    "1111010011111011",
    "1111011001010011",
    "1111011110000101",
    "1111100001111001",
    "1111100100100100",
    "1111100110001110",
    "1111100111011010",
    "1111101000110101",
    "1111101011000001",
    "1111101110001101",
    "1111110010001110",
    "1111110110100010",
    "1111111010100110",
    "1111111110000100",
    "1111111111000110",
    "1111111100101111",
    "1111111010100011",
    "1111111000011001",
    "1111110110010101",
    "1111110100101010",
    "1111110011101100",
    "1111110011101010",
    "1111110100101010",
    "1111110110100110",
    "1111111001010101",
    "1111111100100011",
    "1111111111110010",
    "1111111101101001",
    "1111111100101000",
    "1111111101110100",
    "1111111110011010",
    "1111111000011011",
    "1111110001000000",
    "1111101001001101",
    "1111100010000101",
    "1111011100001110",
    "1111010111101000",
    "1111010011111011",
    "1111010000011100",
    "1111001100110010",
    "1111001000110000",
    "1111000100110111",
    "1111000001110100",
    "1111000000011001",
    "1111000000111101",
    "1111000011011010",
    "1111000111000110",
    "1111001011000110",
    "1111001110100110",
    "1111010001000010",
    "1111010010010100",
    "1111010010110001",
    "1111010010111011",
    "1111010011010010",
    "1111010100001110",
    "1111010110000000",
    "1111011000100010",
    "1111011011101101",
    "1111011111010001",
    "1111100011000000",
    "1111100111000011",
    "1111101100011001",
    "1111110101000000",
    "1111111101000111",
    "1111101001000000",
    "1111001111010100",
    "1110110010100111",
    "1110010110101000",
    "1101111111010110",
    "1101101111011111",
    "1101100111101101",
    "1101100110101010",
    "1101101001101011",
    "1101101110000100",
    "1101110001111000",
    "1101110100010010",
    "1101110101100000",
    "1101110110010101",
    "1101110111100010",
    "1101111001100011",
    "1101111100011011",
    "1101111111101011",
    "1110000010111011",
    "1110000101110110",
    "1110001000010011",
    "1110001010001111",
    "1110001011101000",
    "1110001100100000",
    "1110001100111111",
    "1110001101011011",
    "1110001110010001",
    "1110010000010100",
    "1110010100110110",
    "1110011101011110",
    "1110101011001001",
    "1110111101101011",
    "1111010011010101",
    "1111101001010011",
    "1111111100101010",
    "1111110100110111",
    "1111101100001011",
    "1111101000011010",
    "1111100111110000",
    "1111101000010000",
    "1111101000100010",
    "1111101000001000",
    "1111100111001011",
    "1111100110001011",
    "1111100101110010",
    "1111100110100010",
    "1111101000110110",
    "1111101100110111",
    "1111110010101000",
    "1111111001110101",
    "1111111110000100",
    "1111110110000011",
    "1111101111001100",
    "1111101010100101",
    "1111101000111001",
    "1111101010001001",
    "1111101101100101",
    "1111110010000100",
    "1111110110010010",
    "1111111001000010",
    "1111111001100101",
    "1111110111110010",
    "1111110100001100",
    "1111101111111110",
    "1111101100011100",
    "1111101010110010",
    "1111101011101101",
    "1111101111011100",
    "1111110101101111",
    "1111111110000100",
    "1111111000001111",
    "1111101110001010",
    "1111100100101111",
    "1111011101001111",
    "1111011000101000",
    "1111010111011011",
    "1111011001011101",
    "1111011110000010",
    "1111100100000000",
    "1111101010001000",
    "1111101111010010",
    "1111110010011100",
    "1111110010110100",
    "1111101111110111",
    "1111101001011101",
    "1111011111111111",
    "1111010100011100",
    "1111001000010000",
    "1110111101000101",
    "1110110100011010",
    "1110101111001000",
    "1110101101100000",
    "1110101111000010",
    "1110110010111001",
    "1110111000001000",
    "1110111101101001",
    "1111000010100010",
    "1111000101111011",
    "1111000111000100",
    "1111000101100101",
    "1111000001100001",
    "1110111011101000",
    "1110110101000101",
    "1110101111000100",
    "1110101010101000",
    "1110101000001110",
    "1110100111101101",
    "1110101000101100",
    "1110101010100010",
    "1110101100110101",
    "1110101111011111",
    "1110110010100100",
    "1110110110001110",
    "1110111010100010",
    "1110111111011111",
    "1111000100111100",
    "1111001010100101",
    "1111001111111111",
    "1111010100110011",
    "1111011000110000",
    "1111011011111000",
    "1111011110100011",
    "1111100001010111",
    "1111100100111110",
    "1111101001110010",
    "1111101111101010",
    "1111110110000000",
    "1111111011111001",
    "1111111111100100",
    "1111111101000111",
    "1111111101000001",
    "1111111111001100",
    "1111111100101110",
    "1111110111011010",
    "1111110001100010",
    "1111101011110101",
    "1111100110111011",
    "1111100011010011",
    "1111100001010111",
    "1111100001010000",
    "1111100010111001",
    "1111100110001001",
    "1111101010101110",
    "1111110000011000",
    "1111110110111011",
    "1111111110001111",
    "1111111001111011",
    "1111110010001011",
    "1111101011001111",
    "1111100101111001",
    "1111100010110110",
    "1111100010011001",
    "1111100100100000",
    "1111101000110101",
    "1111101110111010",
    "1111110110010100",
    "1111111110101001",
    "1111111000100010",
    "1111101111111001",
    "1111101000000010",
    "1111100001011100",
    "1111011100010011",
    "1111011000011110",
    "1111010101100101",
    "1111010011001000",
    "1111010000111000",
    "1111001110110110",
    "1111001101100000",
    "1111001101010110",
    "1111001110111000",
    "1111010010010000",
    "1111010111000100",
    "1111011100010111",
    "1111100000111101",
    "1111100011101100",
    "1111100011111001",
    "1111100001011111",
    "1111011101001010",
    "1111011000001000",
    "1111010011110100",
    "1111010001100001",
    "1111010010000011",
    "1111010101100010",
    "1111011011011101",
    "1111100010110011",
    "1111101010100011",
    "1111110001110110",
    "1111111000001111",
    "1111111101101010",
    "1111111101101011",
    "1111111001100100",
    "1111110101110111",
    "1111110010100101",
    "1111101111111000",
    "1111101101111110",
    "1111101101001001",
    "1111101101101100",
    "1111101111101101",
    "1111110011001011",
    "1111110111101111",
    "1111111100110100",
    "1111111110010001",
    "1111111010010001",
    "1111110111101001",
    "1111110110100000",
    "1111110110110100",
    "1111111000010101",
    "1111111010111100",
    "1111111110100100",
    "1111111100101010",
    "1111110110110001",
    "1111101111110101",
    "1111101000001000",
    "1111100000010001",
    "1111011000111110",
    "1111010011000011",
    "1111001111000101",
    "1111001101100001",
    "1111001110011011",
    "1111010001101100",
    "1111010110111110",
    "1111011101011110",
    "1111100100011000",
    "1111101010100111",
    "1111101111010101",
    "1111110010000000",
    "1111110010101001",
    "1111110001101011",
    "1111101111111110",
    "1111101110011110",
    "1111101110000001",
    "1111101111001101",
    "1111110010001011",
    "1111110110101100",
    "1111111100000110",
    "1111111110010111",
    "1111111001100100",
    "1111110101111001",
    "1111110011010011",
    "1111110001010000",
    "1111101110111111",
    "1111101011110100",
    "1111100111011101",
    "1111100010001000",
    "1111011100100110",
    "1111010111111010",
    "1111010101000101",
    "1111010100111001",
    "1111010111110010",
    "1111011101110010",
    "1111100110101011",
    "1111110010000110",
    "1111111111011011",
    "1111110010001101",
    "1111100011111100",
    "1111010110110110",
    "1111001011110000",
    "1111000011001011",
    "1110111101000101",
    "1110111001001110",
    "1110110111000110",
    "1110110110010110",
    "1110110110110001",
    "1110111000001100",
    "1110111010100101",
    "1110111101110101",
    "1111000001111011",
    "1111000110101100",
    "1111001011111010",
    "1111010001010100",
    "1111010110010110",
    "1111011010100110",
    "1111011101101101",
    "1111011111100100",
    "1111100000011110",
    "1111100000111011",
    "1111100001100111",
    "1111100010111110",
    "1111100101001011",
    "1111100111111100",
    "1111101010101100",
    "1111101100110100",
    "1111101101110110",
    "1111101101101101",
    "1111101100110000",
    "1111101011101001",
    "1111101011001001",
    "1111101011110101",
    "1111101101110101",
    "1111110000110001",
    "1111110011111010",
    "1111110110011010",
    "1111110111100111",
    "1111110111011000",
    "1111110110001100",
    "1111110100111100",
    "1111110100100110",
    "1111110101110101",
    "1111111000110001",
    "1111111100111100",
    "1111111110100001",
    "1111111010100011",
    "1111110111101011",
    "1111110101101100",
    "1111110011110111",
    "1111110001001000",
    "1111101100100110",
    "1111100101110110",
    "1111011101001100",
    "1111010011011000",
    "1111001001100011",
    "1111000000110000",
    "1110111001111010",
    "1110110101011101",
    "1110110011011111",
    "1110110011101010",
    "1110110101011011",
    "1110111000001000",
    "1110111011000111",
    "1110111101111010",
    "1111000000010100",
    "1111000010010101",
    "1111000100001101",
    "1111000110001000",
    "1111001000010001",
    "1111001010101101",
    "1111001101010110",
    "1111010000000101",
    "1111010010101110",
    "1111010101010010",
    "1111010111110010",
    "1111011010011011",
    "1111011101011100",
    "1111100001100010",
    "1111101000100101",
    "1111110101000101",
    "1111110111000010",
    "1111011011110010",
    "1110111011101101",
    "1110011011010011",
    "1101111111101000",
    "1101101100111010",
    "1101100100110011",
    "1101100101111110",
    "1101101100111101",
    "1101110101101111",
    "1101111101000101",
    "1110000001100110",
    "1110000011010010",
    "1110000011010111",
    "1110000011001011",
    "1110000011101001",
    "1110000100111001",
    "1110000110100101",
    "1110001000000100",
    "1110001000111111",
    "1110001001011011",
    "1110001001101011",
    "1110001010000010",
    "1110001010100010",
    "1110001011000100",
    "1110001011110101",
    "1110001101001001",
    "1110001111110001",
    "1110010101000011",
    "1110011110011111",
    "1110101101001001",
    "1111000000111000",
    "1111010111111100",
    "1111101111010100",
    "1111111100011001",
    "1111101110000011",
    "1111100110110010",
    "1111100101110110",
    "1111101001000100",
    "1111101101110101",
    "1111110001111100",
    "1111110100001101",
    "1111110100010101",
    "1111110010101010",
    "1111101111111010",
    "1111101100111101",
    "1111101010100110",
    "1111101001100010",
    "1111101010001111",
    "1111101100111110",
    "1111110001110011",
    "1111111000100001",
    "1111111111010111",
    "1111110110101100",
    "1111101110010100",
    "1111100111000001",
    "1111100001010101",
    "1111011101101001",
    "1111011100010011",
    "1111011101100001",
    "1111100001011110",
    "1111101000000001",
    "1111110000101001",
    "1111111010011001",
    "1111111100000010",
    "1111110100000100",
    "1111101110101101",
    "1111101100010101",
    "1111101100100110",
    "1111101110101001",
    "1111110001010111",
    "1111110011110000",
    "1111110101001110",
    "1111110101101010",
    "1111110101010111",
    "1111110100110001",
    "1111110100010001",
    "1111110100000011",
    "1111110100000101",
    "1111110100001010",
    "1111110011111110",
    "1111110011001000",
    "1111110001001110",
    "1111101110000011",
    "1111101001100110",
    "1111100100000110",
    "1111011110000000",
    "1111010111111010",
    "1111010010010100",
    "1111001101100000",
    "1111001001011011",
    "1111000101101100",
    "1111000001110001",
    "1110111101001111",
    "1110110111111111",
    "1110110010011010",
    "1110101101010001",
    "1110101001100101",
    "1110101000001110",
    "1110101001101011",
    "1110101101110000",
    "1110110011100100",
    "1110111001101101",
    "1110111110101000",
    "1111000001000000",
    "1111000000001101",
    "1110111100011001",
    "1110110110011011",
    "1110101111101011",
    "1110101001100101",
    "1110100101011011",
    "1110100100001000",
    "1110100110001011",
    "1110101011100011",
    "1110110011101110",
    "1110111101101101",
    "1111001000001110",
    "1111010001111011",
    "1111011001110010",
    "1111011111010001",
    "1111100010011100",
    "1111100011110110",
    "1111100100001101",
    "1111100100001000",
    "1111100011111100",
    "1111100011101100",
    "1111100011001111",
    "1111100010100001",
    "1111100001101001",
    "1111100000111110",
    "1111100000111110",
    "1111100010001010",
    "1111100100110111",
    "1111101001000101",
    "1111101110011110",
    "1111110100010000",
    "1111111001011111",
    "1111111101010010",
    "1111111111000011",
    "1111111110110000",
    "1111111101000001",
    "1111111010110111",
    "1111111001011001",
    "1111111001011100",
    "1111111011010000",
    "1111111110100010",
    "1111111101011100",
    "1111111001101011",
    "1111110110111010",
    "1111110101101111",
    "1111110110011111",
    "1111111001001110",
    "1111111101110001",
    "1111111100001101",
    "1111110101011010",
    "1111101110011110",
    "1111100111111101",
    "1111100010001111",
    "1111011101010111",
    "1111011001001100",
    "1111010101011101",
    "1111010010000011",
    "1111001111000100",
    "1111001100111000",
    "1111001011111100",
    "1111001100101101",
    "1111001111010110",
    "1111010011101111",
    "1111011001100011",
    "1111011111111011",
    "1111100101111001",
    "1111101010010010",
    "1111101100001010",
    "1111101010111000",
    "1111100110100010",
    "1111011111111101",
    "1111011000100010",
    "1111010001111011",
    "1111001101101110",
    "1111001100110101",
    "1111001111100001",
    "1111010101010101",
    "1111011101011100",
    "1111100111000010",
    "1111110001011000",
    "1111111100000111",
    "1111111001000000",
    "1111101110011011",
    "1111100100101001",
    "1111011100100000",
    "1111010110110111",
    "1111010100100010",
    "1111010101111011",
    "1111011011000110",
    "1111100011011111",
    "1111101110000000",
    "1111111001001001",
    "1111111100101110",
    "1111110101000001",
    "1111110000100011",
    "1111101111011011",
    "1111110001000110",
    "1111110100101011",
    "1111111001001011",
    "1111111101111000",
    "1111111101011100",
    "1111111000110001",
    "1111110011101110",
    "1111101101111010",
    "1111100111000101",
    "1111011111010010",
    "1111010110111001",
    "1111001110101001",
    "1111000111011000",
    "1111000001111000",
    "1110111110101011",
    "1110111110000101",
    "1111000000000000",
    "1111000011111011",
    "1111001001000111",
    "1111001110110001",
    "1111010100000101",
    "1111011000100011",
    "1111011011111111",
    "1111011110011110",
    "1111100000010100",
    "1111100001111011",
    "1111100011110001",
    "1111100110001000",
    "1111101001001111",
    "1111101101000101",
    "1111110001011010",
    "1111110101111000",
    "1111111010001000",
    "1111111110000001",
    "1111111110001101",
    "1111111010000110",
    "1111110100111110",
    "1111101110011101",
    "1111100110101001",
    "1111011110010010",
    "1111010110100010",
    "1111010000101001",
    "1111001101101000",
    "1111001101111101",
    "1111010001011111",
    "1111010111101100",
    "1111011111110011",
    "1111101001001001",
    "1111110011000011",
    "1111111100111110",
    "1111111001100010",
    "1111110001000000",
    "1111101001101111",
    "1111100011111110",
    "1111011111110000",
    "1111011100111111",
    "1111011011011001",
    "1111011010100000",
    "1111011001110100",
    "1111011000110010",
    "1111010110110111",
    "1111010011110001",
    "1111001111011110",
    "1111001010011000",
    "1111000101001110",
    "1111000000111001",
    "1110111110001100",
    "1110111101101000",
    "1110111111011100",
    "1111000011100111",
    "1111001001110101",
    "1111010001101011",
    "1111011010010011",
    "1111100010110001",
    "1111101001111111",
    "1111101110111110",
    "1111110001001010",
    "1111110000100111",
    "1111101110001011",
    "1111101011000011",
    "1111101000101100",
    "1111101000001011",
    "1111101010000100",
    "1111101110001000",
    "1111110011100010",
    "1111111001000110",
    "1111111101100110",
    "1111111111111011",
    "1111111111111100",
    "1111111101011011",
    "1111111001001100",
    "1111110100010101",
    "1111101111111100",
    "1111101100111101",
    "1111101011110000",
    "1111101100001100",
    "1111101101110000",
    "1111101111110100",
    "1111110001111101",
    "1111110100001111",
    "1111110111000101",
    "1111111011001001",
    "1111111111000101",
    "1111110111100011",
    "1111101110100111",
    "1111100100111100",
    "1111011011011001",
    "1111010010100110",
    "1111001010111000",
    "1111000100011000",
    "1110111111000111",
    "1110111011010001",
    "1110111001001110",
    "1110111001010001",
    "1110111011011101",
    "1110111111011010",
    "1111000100011000",
    "1111001001010110",
    "1111001101011001",
    "1111010000000010",
    "1111010001001010",
    "1111010001001111",
    "1111010000110000",
    "1111010000010101",
    "1111010000010101",
    "1111010000111101",
    "1111010010001010",
    "1111010011111001",
    "1111010110000110",
    "1111011000101111",
    "1111011011110000",
    "1111011111001100",
    "1111100011011111",
    "1111101010010001",
    "1111110101111011",
    "1111110111011111",
    "1111011101101101",
    "1110111110110000",
    "1110011110101101",
    "1110000010011100",
    "1101101110010010",
    "1101100100010011",
    "1101100011101111",
    "1101101001110010",
    "1101110010101011",
    "1101111011010110",
    "1110000010000110",
    "1110000110101010",
    "1110001001100011",
    "1110001011101111",
    "1110001101101000",
    "1110001111001101",
    "1110010000000111",
    "1110001111110110",
    "1110001110011011",
    "1110001100001100",
    "1110001001111010",
    "1110001000001001",
    "1110000111001001",
    "1110000110111110",
    "1110000111101101",
    "1110001001100101",
    "1110001100111000",
    "1110010010000000",
    "1110011001010110",
    "1110100011011010",
    "1110110000011100",
    "1111000000010111",
    "1111010010101011",
    "1111100110100001",
    "1111111010110110",
    "1111110001100111",
    "1111100000010001",
    "1111010010010101",
    "1111001000111110",
    "1111000100110110",
    "1111000110000011",
    "1111001100000010",
    "1111010101110001",
    "1111100001111001",
    "1111101111001001",
    "1111111100001111",
    "1111110111111110",
    "1111101110101001",
    "1111101000100111",
    "1111100110010011",
    "1111100111100001",
    "1111101011011001",
    "1111110000101111",
    "1111110110100100",
    "1111111100001000",
    "1111111110111001",
    "1111111010110001",
    "1111110111100111",
    "1111110101110000",
    "1111110101110000",
    "1111111000000111",
    "1111111100110111",
    "1111111100011011",
    "1111110101000001",
    "1111101110010100",
    "1111101001110001",
    "1111101000011010",
    "1111101010110010",
    "1111110000110100",
    "1111111001111001",
    "1111111011000001",
    "1111101111011100",
    "1111100100110111",
    "1111011100101101",
    "1111010111101101",
    "1111010101111100",
    "1111010110101100",
    "1111011000101101",
    "1111011010101111",
    "1111011011111010",
    "1111011011110101",
    "1111011010100011",
    "1111011000010011",
    "1111010101010101",
    "1111010001110100",
    "1111001101110011",
    "1111001001010101",
    "1111000100011101",
    "1110111111100001",
    "1110111010110100",
    "1110110110101010",
    "1110110011010111",
    "1110110001000111",
    "1110101111111011",
    "1110101111111010",
    "1110110000111000",
    "1110110010101011",
    "1110110100111001",
    "1110110111000011",
    "1110111000100010",
    "1110111000111001",
    "1110110111111001",
    "1110110101100010",
    "1110110010000110",
    "1110101110000100",
    "1110101010000001",
    "1110100110101010",
    "1110100100100100",
    "1110100100001010",
    "1110100101100111",
    "1110101000111100",
    "1110101101111010",
    "1110110100001101",
    "1110111011011101",
    "1111000011010010",
    "1111001011010100",
    "1111010011001011",
    "1111011010011110",
    "1111100000110110",
    "1111100110000011",
    "1111101001111111",
    "1111101100101001",
    "1111101110000011",
    "1111101110010101",
    "1111101101100101",
    "1111101011111101",
    "1111101001101001",
    "1111100110111110",
    "1111100100010101",
    "1111100010001101",
    "1111100000111110",
    "1111100000110110",
    "1111100001110100",
    "1111100011101001",
    "1111100101111100",
    "1111101000100101",
    "1111101011100001",
    "1111101111001000",
    "1111110011111001",
    "1111111010001100",
    "1111111101111011",
    "1111110101001001",
    "1111101100100010",
    "1111100101011101",
    "1111100001000111",
    "1111100000001010",
    "1111100010100111",
    "1111100111110011",
    "1111101110101001",
    "1111110110000100",
    "1111111101001001",
    "1111111100100000",
    "1111110110111111",
    "1111110010000110",
    "1111101101100110",
    "1111101001011101",
    "1111100101111001",
    "1111100011010011",
    "1111100010001101",
    "1111100010111000",
    "1111100101001110",
    "1111101000110101",
    "1111101100110100",
    "1111110000010001",
    "1111110010010000",
    "1111110010001000",
    "1111101111011111",
    "1111101010010010",
    "1111100010111011",
    "1111011010001100",
    "1111010001001101",
    "1111001001010011",
    "1111000011110011",
    "1111000001101100",
    "1111000011100001",
    "1111001001000110",
    "1111010001101100",
    "1111011100001100",
    "1111100111010000",
    "1111110001110001",
    "1111111010110101",
    "1111111110000011",
    "1111111001001100",
    "1111110110100001",
    "1111110101110011",
    "1111110110101010",
    "1111111000110010",
    "1111111011111010",
    "1111111111110110",
    "1111111011100110",
    "1111110110110111",
    "1111110010100010",
    "1111101111011001",
    "1111101110010001",
    "1111101111100010",
    "1111110011000010",
    "1111110111111110",
    "1111111101001010",
    "1111111110011111",
    "1111111011101101",
    "1111111010011101",
    "1111111010001001",
    "1111111001111010",
    "1111111000111011",
    "1111110110101111",
    "1111110011010011",
    "1111101110111010",
    "1111101010000110",
    "1111100101011000",
    "1111100001010000",
    "1111011110001001",
    "1111011100010001",
    "1111011011110010",
    "1111011100100110",
    "1111011110010111",
    "1111100000100110",
    "1111100010101001",
    "1111100100000000",
    "1111100100010101",
    "1111100011100100",
    "1111100001111110",
    "1111100000000011",
    "1111011110011011",
    "1111011101101101",
    "1111011110011111",
    "1111100000111110",
    "1111100101000110",
    "1111101010010110",
    "1111110000000011",
    "1111110101100010",
    "1111111010010111",
    "1111111110100000",
    "1111111101101100",
    "1111111001110010",
    "1111110101011101",
    "1111110000101100",
    "1111101011111000",
    "1111100111101101",
    "1111100100110100",
    "1111100011100110",
    "1111100011111110",
    "1111100101100100",
    "1111100111101111",
    "1111101001111001",
    "1111101011110000",
    "1111101101011010",
    "1111101111010110",
    "1111110010010001",
    "1111110110111111",
    "1111111110000010",
    "1111111000011111",
    "1111101101001101",
    "1111100001001000",
    "1111010101101001",
    "1111001011111000",
    "1111000100101111",
    "1111000000011001",
    "1110111110011111",
    "1110111110011001",
    "1110111111011100",
    "1111000001001101",
    "1111000011100100",
    "1111000110100010",
    "1111001010000010",
    "1111001101111000",
    "1111010001101100",
    "1111010100111110",
    "1111010111011101",
    "1111011000111111",
    "1111011001101111",
    "1111011001110111",
    "1111011001100011",
    "1111011000111001",
    "1111010111111111",
    "1111010111000001",
    "1111010110010011",
    "1111010110010101",
    "1111010111100000",
    "1111011010000001",
    "1111011101101101",
    "1111100010000110",
    "1111100110011111",
    "1111101010001010",
    "1111101100101000",
    "1111101101101111",
    "1111101101101100",
    "1111101100111100",
    "1111101100000010",
    "1111101011011100",
    "1111101011010101",
    "1111101011101000",
    "1111101011111001",
    "1111101011100000",
    "1111101001111110",
    "1111100111001100",
    "1111100011100001",
    "1111011111110110",
    "1111011101011011",
    "1111011101011110",
    "1111100001000010",
    "1111101000100010",
    "1111110011110000",
    "1111111110010000",
    "1111101111001010",
    "1111100000101011",
    "1111010100010111",
    "1111001011000111",
    "1111000101000011",
    "1111000001100111",
    "1110111111111101",
    "1110111111001111",
    "1110111111000101",
    "1110111111011001",
    "1111000000010001",
    "1111000001110011",
    "1111000011110011",
    "1111000101110111",
    "1111000111100101",
    "1111001000100101",
    "1111001000110010",
    "1111001000010110",
    "1111000111100111",
    "1111000110111001",
    "1111000110011011",
    "1111000110010110",
    "1111000110101000",
    "1111000111010011",
    "1111001000011101",
    "1111001010001111",
    "1111001100110111",
    "1111010000010101",
    "1111010100110001",
    "1111011010011101",
    "1111100010101110",
    "1111101111100111",
    "1111111101001001",
    "1111100011010101",
    "1111000100110100",
    "1110100101011101",
    "1110001001110101",
    "1101110110001001",
    "1101101100011011",
    "1101101100000010",
    "1101110010001011",
    "1101111011000001",
    "1110000011001000",
    "1110001000100101",
    "1110001010110101",
    "1110001010101000",
    "1110001001001110",
    "1110000111101100",
    "1110000110100111",
    "1110000110001001",
    "1110000110000110",
    "1110000110010101",
    "1110000110111001",
    "1110000111110111",
    "1110001001001011",
    "1110001010100110",
    "1110001011110111",
    "1110001100111010",
    "1110001110001010",
    "1110010000010001",
    "1110010100100100",
    "1110011100111000",
    "1110101011000100",
    "1110111111111000",
    "1111011010001001",
    "1111110110110000",
    "1111101110011111",
    "1111011001110101",
    "1111001110000101",
    "1111001011110101",
    "1111010001011100",
    "1111011011101111",
    "1111100111010000",
    "1111110001010110",
    "1111111000100101",
    "1111111100101000",
    "1111111110001011",
    "1111111110010111",
    "1111111110010100",
    "1111111110110011",
    "1111111111110011",
    "1111111101101001",
    "1111111010110111",
    "1111110111101010",
    "1111110100001101",
    "1111110000110011",
    "1111101101111000",
    "1111101011110100",
    "1111101010110010",
    "1111101010111001",
    "1111101100001100",
    "1111101110101101",
    "1111110010010110",
    "1111110110110101",
    "1111111011101101",
    "1111111111100000",
    "1111111011011001",
    "1111111000010011",
    "1111110110011010",
    "1111110101100100",
    "1111110101011001",
    "1111110101011110",
    "1111110101100001",
    "1111110101010100",
    "1111110100110111",
    "1111110100001111",
    "1111110011100100",
    "1111110010110110",
    "1111110010000101",
    "1111110001000110",
    "1111101111111010",
    "1111101110100100",
    "1111101101001101",
    "1111101011110100",
    "1111101010001101",
    "1111100111111110",
    "1111100100101001",
    "1111011111111010",
    "1111011001101101",
    "1111010010011010",
    "1111001010101101",
    "1111000011011101",
    "1110111101100110",
    "1110111001101101",
    "1110110111111010",
    "1110110111110111",
    "1110111000101111",
    "1110111001100010",
    "1110111001010000",
    "1110110111011011",
    "1110110100001011",
    "1110110000001100",
    "1110101100010001",
    "1110101001001100",
    "1110100111010000",
    "1110100110010101",
    "1110100101111110",
    "1110100101110100",
    "1110100101110001",
    "1110100110000100",
    "1110100111001101",
    "1110101001100101",
    "1110101101011100",
    "1110110010101110",
    "1110111001000100",
    "1110111111111101",
    "1111000110111001",
    "1111001101010110",
    "1111010010111000",
    "1111010111001101",
    "1111011010001001",
    "1111011011101000",
    "1111011011110010",
    "1111011010110010",
    "1111011000111111",
    "1111010110110111",
    "1111010100111110",
    "1111010011110100",
    "1111010011110110",
    "1111010101001101",
    "1111010111101010",
    "1111011010110010",
    "1111011101111010",
    "1111100000100100",
    "1111100010100110",
    "1111100100011000",
    "1111100110101010",
    "1111101010001111",
    "1111101111100011",
    "1111110110011111",
    "1111111110001100",
    "1111111010101011",
    "1111110101100101",
    "1111110011100110",
    "1111110101001001",
    "1111111001111000",
    "1111111111000110",
    "1111110111000110",
    "1111101111011010",
    "1111101001001001",
    "1111100100111110",
    "1111100011000101",
    "1111100011010010",
    "1111100100111100",
    "1111100111011000",
    "1111101001110100",
    "1111101011101111",
    "1111101100110101",
    "1111101101000101",
    "1111101100100010",
    "1111101011010100",
    "1111101001100001",
    "1111100111001101",
    "1111100100011010",
    "1111100001001111",
    "1111011101110000",
    "1111011010001100",
    "1111010110101100",
    "1111010011011101",
    "1111010000101001",
    "1111001110011001",
    "1111001100111000",
    "1111001100010011",
    "1111001100110101",
    "1111001110100001",
    "1111010001001100",
    "1111010100100000",
    "1111011000000100",
    "1111011011101000",
    "1111011111001010",
    "1111100011000011",
    "1111100111110101",
    "1111101101111111",
    "1111110101101010",
    "1111111110011001",
    "1111111000101010",
    "1111110000111000",
    "1111101011011100",
    "1111101001001100",
    "1111101010011001",
    "1111101110101000",
    "1111110100111010",
    "1111111011111000",
    "1111111101101101",
    "1111111000111000",
    "1111110110000000",
    "1111110100111010",
    "1111110101000011",
    "1111110101110001",
    "1111110110101011",
    "1111110111101101",
    "1111111001001100",
    "1111111011100000",
    "1111111111000010",
    "1111111100001010",
    "1111110110011001",
    "1111110000001000",
    "1111101001111001",
    "1111100100001101",
    "1111011111011001",
    "1111011011101010",
    "1111011000111100",
    "1111010111000011",
    "1111010101101100",
    "1111010100011010",
    "1111010010110100",
    "1111010000100111",
    "1111001101110011",
    "1111001010100110",
    "1111000111100000",
    "1111000101001000",
    "1111000100000011",
    "1111000100110011",
    "1111000111100101",
    "1111001100010100",
    "1111010010100111",
    "1111011001101000",
    "1111100000011001",
    "1111100110000011",
    "1111101001111100",
    "1111101100000100",
    "1111101100111101",
    "1111101101100101",
    "1111101110111111",
    "1111110001111010",
    "1111110110100110",
    "1111111100110011",
    "1111111100000010",
    "1111110100101100",
    "1111101101110110",
    "1111100111111010",
    "1111100011001011",
    "1111011111110001",
    "1111011101111000",
    "1111011101101000",
    "1111011111000111",
    "1111100010011111",
    "1111100111101101",
    "1111101110100111",
    "1111110110110001",
    "1111111111011110",
    "1111111000001011",
    "1111110001000110",
    "1111101011111101",
    "1111101001000001",
    "1111100111111111",
    "1111101000001001",
    "1111101000010011",
    "1111100111010000",
    "1111100100000110",
    "1111011110100110",
    "1111010111010000",
    "1111001111001100",
    "1111000111110101",
    "1111000010010101",
    "1110111111011001",
    "1110111111000010",
    "1111000000110101",
    "1111000100000001",
    "1111000111111001",
    "1111001011110000",
    "1111001111000111",
    "1111010001101001",
    "1111010011001111",
    "1111010100001010",
    "1111010100110110",
    "1111010110000000",
    "1111011000001000",
    "1111011011100011",
    "1111100000010001",
    "1111100101110110",
    "1111101011101101",
    "1111110001001000",
    "1111110101100010",
    "1111111000100011",
    "1111111010000011",
    "1111111010001001",
    "1111111001000011",
    "1111110111000010",
    "1111110100010011",
    "1111110000111111",
    "1111101101001001",
    "1111101000110011",
    "1111100100000110",
    "1111011111010111",
    "1111011011001010",
    "1111011000010000",
    "1111010111010000",
    "1111011000100111",
    "1111011100010001",
    "1111100001110100",
    "1111101000101001",
    "1111110000000010",
    "1111110111100010",
    "1111111111000001",
    "1111111001011011",
    "1111110001101101",
    "1111101001110011",
    "1111100001111011",
    "1111011010011101",
    "1111010011110110",
    "1111001110011100",
    "1111001010100011",
    "1111001000010011",
    "1111000111101100",
    "1111001000011110",
    "1111001010010011",
    "1111001100100011",
    "1111001110100110",
    "1111001111110110",
    "1111010000000010",
    "1111001111001111",
    "1111001101110101",
    "1111001100011001",
    "1111001011100000",
    "1111001011100001",
    "1111001100100101",
    "1111001110100011",
    "1111010001001000",
    "1111010100000000",
    "1111010110111110",
    "1111011001111100",
    "1111011100111000",
    "1111011111111011",
    "1111100011001011",
    "1111100111010010",
    "1111101110001100",
    "1111111010100110",
    "1111110001011011",
    "1111010101111011",
    "1110110101100010",
    "1110010101000001",
    "1101111001101101",
    "1101100111111010",
    "1101100001010010",
    "1101100100010000",
    "1101101101001100",
    "1101110111101111",
    "1110000000100100",
    "1110000110001101",
    "1110001000100011",
    "1110001000101101",
    "1110000111111100",
    "1110000111000011",
    "1110000110010000",
    "1110000101011011",
    "1110000100010111",
    "1110000011000101",
    "1110000010001000",
    "1110000010000010",
    "1110000011000011",
    "1110000101000001",
    "1110000111100101",
    "1110001010100101",
    "1110001110000010",
    "1110010010001010",
    "1110010111100010",
    "1110011111000111",
    "1110101001110010",
    "1110111000000001",
    "1111001001011000",
    "1111011100100011",
    "1111101111101011",
    "1111111111000100",
    "1111110001001101",
    "1111100111011100",
    "1111100001110001",
    "1111011111110000",
    "1111100000111000",
    "1111100100101100",
    "1111101010101010",
    "1111110010000110",
    "1111111010000111",
    "1111111110001011",
    "1111110111110001",
    "1111110011010110",
    "1111110001011111",
    "1111110010001111",
    "1111110101010000",
    "1111111001101010",
    "1111111110011100",
    "1111111101010100",
    "1111111010010010",
    "1111111000100100",
    "1111111000000010",
    "1111111000010100",
    "1111111000111011",
    "1111111001011111",
    "1111111001111010",
    "1111111010011000",
    "1111111011001100",
    "1111111100100011",
    "1111111110011011",
    "1111111111011000",
    "1111111101010011",
    "1111111011111001",
    "1111111011101010",
    "1111111101000100",
    "1111111111100111",
    "1111111010010111",
    "1111110011010111",
    "1111101011001011",
    "1111100010100100",
    "1111011010011101",
    "1111010011101001",
    "1111001110101101",
    "1111001011110111",
    "1111001011000110",
    "1111001011111111",
    "1111001101110011",
    "1111001111101011",
    "1111010000100111",
    "1111001111111011",
    "1111001101010010",
    "1111001000111001",
    "1111000011010000",
    "1110111101001110",
    "1110110111100111",
    "1110110010110110",
    "1110101111000010",
    "1110101011110101",
    "1110101000110101",
    "1110100101110010",
    "1110100010110001",
    "1110100000001101",
    "1110011110101110",
    "1110011110101110",
    "1110100000001111",
    "1110100010101110",
    "1110100101001101",
    "1110100110101101",
    "1110100110101010",
    "1110100100111011",
    "1110100010000011",
    "1110011111000010",
    "1110011101000111",
    "1110011101010001",
    "1110100000001010",
    "1110100101111011",
    "1110101110001100",
    "1110111000010001",
    "1111000011001101",
    "1111001101101110",
    "1111010110101111",
    "1111011101010010",
    "1111100000110101",
    "1111100001010010",
    "1111011111000101",
    "1111011010111100",
    "1111010101101111",
    "1111010000011110",
    "1111001011111101",
    "1111001000111110",
    "1111000111110111",
    "1111001000101101",
    "1111001011010001",
    "1111001111000010",
    "1111010011100110",
    "1111011000101000",
    "1111011110001001",
    "1111100100010010",
    "1111101011001101",
    "1111110010110001",
    "1111111010011001",
    "1111111110110001",
    "1111111001110000",
    "1111110111001010",
    "1111110111000000",
    "1111111000101101",
    "1111111011010001",
    "1111111101101100",
    "1111111111001100",
    "1111111111100010",
    "1111111110111001",
    "1111111101110101",
    "1111111101000001",
    "1111111100111100",
    "1111111101110000",
    "1111111111011001",
    "1111111110010111",
    "1111111011110110",
    "1111111001001100",
    "1111110110011011",
    "1111110011100010",
    "1111110000100100",
    "1111101101100110",
    "1111101010110011",
    "1111101000010001",
    "1111100101111110",
    "1111100011110001",
    "1111100001011010",
    "1111011110101101",
    "1111011011100101",
    "1111011000000100",
    "1111010100011100",
    "1111010000111101",
    "1111001110000101",
    "1111001100001110",
    "1111001011101011",
    "1111001100101110",
    "1111001111100011",
    "1111010100001000",
    "1111011010011011",
    "1111100010001010",
    "1111101010110101",
    "1111110011101110",
    "1111111100000001",
    "1111111101001001",
    "1111111000100101",
    "1111110110110110",
    "1111111000001000",
    "1111111100010010",
    "1111111101010011",
    "1111110101110001",
    "1111101110011010",
    "1111101000100001",
    "1111100101001101",
    "1111100100111100",
    "1111100111101000",
    "1111101100011111",
    "1111110010010111",
    "1111111000000001",
    "1111111100011101",
    "1111111111000001",
    "1111111111100101",
    "1111111110011110",
    "1111111100010010",
    "1111111001110011",
    "1111110111110001",
    "1111110110110111",
    "1111110111011110",
    "1111111001110001",
    "1111111101100100",
    "1111111101011011",
    "1111110111110001",
    "1111110001110011",
    "1111101011111011",
    "1111100110011010",
    "1111100001011100",
    "1111011101001110",
    "1111011001110101",
    "1111010111011011",
    "1111010110001001",
    "1111010110000000",
    "1111010110110001",
    "1111011000000110",
    "1111011001100000",
    "1111011010100010",
    "1111011010111101",
    "1111011011000001",
    "1111011011001001",
    "1111011100000001",
    "1111011110000101",
    "1111100001011100",
    "1111100101110100",
    "1111101010110010",
    "1111101111110011",
    "1111110100011101",
    "1111111000100010",
    "1111111100000000",
    "1111111111000010",
    "1111111110001001",
    "1111111011010110",
    "1111111000010100",
    "1111110100111011",
    "1111110001001100",
    "1111101101010001",
    "1111101001100110",
    "1111100110101001",
    "1111100101000000",
    "1111100101000101",
    "1111100111001111",
    "1111101011100110",
    "1111110010000011",
    "1111111010100001",
    "1111111011001011",
    "1111101111100110",
    "1111100011100110",
    "1111011000011010",
    "1111001111010111",
    "1111001001010011",
    "1111000110011010",
    "1111000110000011",
    "1111000111001000",
    "1111001000100011",
    "1111001001101111",
    "1111001010100010",
    "1111001011001110",
    "1111001100000101",
    "1111001101010010",
    "1111001110101110",
    "1111010000000101",
    "1111010000111101",
    "1111010001000011",
    "1111010000001111",
    "1111001110101001",
    "1111001100101011",
    "1111001010111101",
    "1111001010001001",
    "1111001010101101",
    "1111001100101011",
    "1111001111101100",
    "1111010011000001",
    "1111010101111110",
    "1111010111111010",
    "1111011000101111",
    "1111011000101010",
    "1111011000000110",
    "1111010111100010",
    "1111010111010101",
    "1111010111100011",
    "1111011000001001",
    "1111011000111100",
    "1111011001101011",
    "1111011010001111",
    "1111011010011001",
    "1111011010000111",
    "1111011001010110",
    "1111011000010000",
    "1111010111000110",
    "1111010110010000",
    "1111010110001001",
    "1111010111001011",
    "1111011001100011",
    "1111011101011001",
    "1111100010110001",
    "1111101001101110",
    "1111110010001111",
    "1111111100001001",
    "1111111000111000",
    "1111101101011100",
    "1111100010010101",
    "1111011000010011",
    "1111010000000010",
    "1111001001110111",
    "1111000101110110",
    "1111000011101010",
    "1111000010110110",
    "1111000010110100",
    "1111000011000101",
    "1111000011010000",
    "1111000011010000",
    "1111000011001011",
    "1111000011001010",
    "1111000011010000",
    "1111000011011111",
    "1111000011110100",
    "1111000100000101",
    "1111000100001110",
    "1111000100010010",
    "1111000100010011",
    "1111000100011111",
    "1111000101000011",
    "1111000110001101",
    "1111001000001000",
    "1111001010111100",
    "1111001110100110",
    "1111010010111011",
    "1111010111100101",
    "1111011100010100",
    "1111100000110110",
    "1111100101010101",
    "1111101010101101",
    "1111110010101011",
    "1111111111000010",
    "1111101111000011",
    "1111010111111100",
    "1110111101101001",
    "1110100011011101",
    "1110001100111111",
    "1101111101000100",
    "1101110100101111",
    "1101110011001111",
    "1101110110011011",
    "1101111011101011",
    "1110000000101110",
    "1110000100010010",
    "1110000110000001",
    "1110000110011000",
    "1110000110000011",
    "1110000101100111",
    "1110000101010010",
    "1110000101000011",
    "1110000100101111",
    "1110000100010010",
    "1110000011111000",
    "1110000011110011",
    "1110000100010000",
    "1110000101011111",
    "1110000111100011",
    "1110001010101101",
    "1110001111000100",
    "1110010101000011",
    "1110011101010010",
    "1110101000011000",
    "1110110110110010",
    "1111001000010101",
    "1111011100001100",
    "1111110000110111",
    "1111111011100100",
    "1111101011000100",
    "1111011111001000",
    "1111011000100111",
    "1111010111110001",
    "1111011100000101",
    "1111100100101010",
    "1111110000000001",
    "1111111100011111",
    "1111110111100111",
    "1111101101101110",
    "1111100110101111",
    "1111100010111001",
    "1111100001111011",
    "1111100011001000",
    "1111100101101010",
    "1111101000110000",
    "1111101011110111",
    "1111101110101110",
    "1111110001010111",
    "1111110011111110",
    "1111110110100110",
    "1111111001001101",
    "1111111011101010",
    "1111111101110000",
    "1111111111001111",
    "1111111111111100",
    "1111111111111101",
    "1111111111000110",
    "1111111101011111",
    "1111111011011100",
    "1111111001010011",
    "1111110111100110",
    "1111110110111000",
    "1111110111100011",
    "1111111001110101",
    "1111111101100110",
    "1111111101100110",
    "1111111000011011",
    "1111110011100011",
    "1111101111011101",
    "1111101100010110",
    "1111101010000110",
    "1111101000010111",
    "1111100110110001",
    "1111100101000001",
    "1111100010111101",
    "1111100000011110",
    "1111011101100100",
    "1111011010010001",
    "1111010110100100",
    "1111010010100001",
    "1111001110010010",
    "1111001001111100",
    "1111000101101001",
    "1111000001011110",
    "1110111101100100",
    "1110111010000001",
    "1110110110110001",
    "1110110011101110",
    "1110110000100100",
    "1110101101000010",
    "1110101000111010",
    "1110100100001010",
    "1110011111000100",
    "1110011010001110",
    "1110010110011011",
    "1110010100011000",
    "1110010100101100",
    "1110010111100101",
    "1110011100111111",
    "1110100100011101",
    "1110101101001110",
    "1110110110010011",
    "1110111110100110",
    "1111000101000110",
    "1111001000111110",
    "1111001001111001",
    "1111000111111111",
    "1111000011111011",
    "1110111110100001",
    "1110111000110111",
    "1110110100000011",
    "1110110001000010",
    "1110110000011100",
    "1110110010100111",
    "1110110111011011",
    "1110111110010100",
    "1111000110100101",
    "1111001111010010",
    "1111010111101010",
    "1111011111000010",
    "1111100101000110",
    "1111101001110010",
    "1111101101010101",
    "1111101111111111",
    "1111110010000010",
    "1111110011100110",
    "1111110100101101",
    "1111110101001111",
    "1111110101001001",
    "1111110100100001"
    );
begin
    
    --clk generator
    clk_gen:process(clk)
    begin
        clk <= not clk after half_period;
    end process;
   
    
    --control stimulus generator
    reset <= '0', '1' after 5ns;
    on_in_s <= '0', '1' after 25ns;
    
    write_output: process(on_in_s, out_valid)
    --declare files/variabbles used for storing output and loading input
    file output_file     : text is out "C:\Users\user\Desktop\text_io_output.txt";
    variable output_line : line;
    variable input_counter: integer := 104590; --hardcoded number of inputs from AUDIO array abve
    begin  
        if out_valid'event then
            if out_valid = '1' then            
                --write new output value to txt file
                write(output_line, std_logic_vector(output_out_s), left, 16);
                writeline (output_file, output_line);
                
                --load new input value
                input_in_s <= AUDIO(input_counter); --load value
                input_counter := input_counter - 1; --decrement counter
            else
            --new input value loaded         
            end if;
        end if;
    end process;
    
    DUT: entity work.phaser_datapath(Behavioral)
                 port map (input_in => input_in_s,
                           on_in => on_in_s,
                           reset => reset,
                           clk => clk,
                           out_valid => out_valid,
                           output_out => output_out_s
                 );
                 

end Behavioral;
